* NGSPICE file created from top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

.subckt top A1[0] A1[1] A1[2] A1[3] A1[4] A2[0] A2[1] A2[2] A2[3] A2[4] A3[0] A3[1]
+ A3[2] A3[3] A3[4] VGND VPWR WD3[0] WD3[10] WD3[11] WD3[12] WD3[13] WD3[14] WD3[15]
+ WD3[16] WD3[17] WD3[18] WD3[19] WD3[1] WD3[20] WD3[21] WD3[22] WD3[23] WD3[24] WD3[25]
+ WD3[26] WD3[27] WD3[28] WD3[29] WD3[2] WD3[30] WD3[31] WD3[3] WD3[4] WD3[5] WD3[6]
+ WD3[7] WD3[8] WD3[9] WE3 alu_out[0] alu_out[10] alu_out[11] alu_out[12] alu_out[13]
+ alu_out[14] alu_out[15] alu_out[16] alu_out[17] alu_out[18] alu_out[19] alu_out[1]
+ alu_out[20] alu_out[21] alu_out[22] alu_out[23] alu_out[24] alu_out[25] alu_out[26]
+ alu_out[27] alu_out[28] alu_out[29] alu_out[2] alu_out[30] alu_out[31] alu_out[3]
+ alu_out[4] alu_out[5] alu_out[6] alu_out[7] alu_out[8] alu_out[9] clk opcode[0]
+ opcode[1]
XANTENNA__6626__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4935__A _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5512__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7963_ net893 _3448_ _3938_ VGND VGND VPWR VPWR _3948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6914_ _3375_ VGND VGND VPWR VPWR _3376_ sky130_fd_sc_hd__buf_4
X_7894_ _3911_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__clkbuf_1
X_6845_ _3091_ _3302_ VGND VGND VPWR VPWR _3339_ sky130_fd_sc_hd__nor2_4
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5766__A _2323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6361__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9564_ clknet_leaf_16_clk _0724_ VGND VGND VPWR VPWR rf.registers\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6776_ net13 net12 net11 VGND VGND VPWR VPWR _3302_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_102_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8515_ _4240_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_99_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5727_ _2062_ _2479_ VGND VGND VPWR VPWR _2480_ sky130_fd_sc_hd__nor2_1
X_9495_ clknet_leaf_33_clk _0655_ VGND VGND VPWR VPWR rf.registers\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7342__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8446_ _3003_ _3411_ VGND VGND VPWR VPWR _4204_ sky130_fd_sc_hd__nor2_4
X_5658_ _2410_ _2412_ _2097_ VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8288__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4609_ _1254_ _1364_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__nor2_1
X_8377_ _4167_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5589_ _1799_ _2141_ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold340 rf.registers\[0\]\[21\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
X_7328_ _3611_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
Xhold351 rf.registers\[22\]\[18\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 rf.registers\[6\]\[18\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 rf.registers\[23\]\[3\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold384 rf.registers\[12\]\[19\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7645__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7259_ _3060_ net964 _3566_ VGND VGND VPWR VPWR _3575_ sky130_fd_sc_hd__mux2_1
Xhold395 rf.registers\[11\]\[23\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1040 rf.registers\[2\]\[6\] VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 rf.registers\[30\]\[29\] VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7221__A _3554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1062 rf.registers\[13\]\[29\] VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4306__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5503__S0 _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7367__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer7 net1167 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4739__B _1480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4545__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output56_A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8061__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4960_ _1655_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__buf_4
X_4891_ rf.registers\[28\]\[0\] rf.registers\[29\]\[0\] rf.registers\[30\]\[0\] rf.registers\[31\]\[0\]
+ net1 net2 VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6630_ _3079_ net996 _3217_ VGND VGND VPWR VPWR _3225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6561_ _3187_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8300_ _3009_ net338 _4119_ VGND VGND VPWR VPWR _4127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5512_ rf.registers\[0\]\[6\] rf.registers\[1\]\[6\] rf.registers\[2\]\[6\] rf.registers\[3\]\[6\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2268_ sky130_fd_sc_hd__mux4_1
X_9280_ clknet_leaf_69_clk _0440_ VGND VGND VPWR VPWR rf.registers\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6492_ _3149_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8231_ _4090_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__clkbuf_1
X_5443_ rf.registers\[16\]\[10\] rf.registers\[17\]\[10\] rf.registers\[18\]\[10\]
+ rf.registers\[19\]\[10\] _2050_ _2052_ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4689__B2 _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6210__A _1996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8162_ net834 _3442_ _4047_ VGND VGND VPWR VPWR _4054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5374_ _2128_ _2129_ _2044_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7113_ net23 VGND VGND VPWR VPWR _3493_ sky130_fd_sc_hd__buf_2
X_4325_ _1079_ _1080_ _1040_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8093_ _4017_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__clkbuf_1
X_7044_ net34 VGND VGND VPWR VPWR _3446_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4536__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4861__B2 _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8052__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8995_ clknet_leaf_67_clk _0155_ VGND VGND VPWR VPWR rf.registers\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7946_ _3939_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4613__A1 _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7877_ _3134_ net689 _3902_ VGND VGND VPWR VPWR _3903_ sky130_fd_sc_hd__mux2_1
XANTENNA__7187__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5496__A _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6828_ _3330_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9547_ clknet_leaf_4_clk _0707_ VGND VGND VPWR VPWR rf.registers\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6759_ _3293_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7915__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6118__A1 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9478_ clknet_leaf_66_clk _0638_ VGND VGND VPWR VPWR rf.registers\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8429_ _4195_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5435__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6120__A _1430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4775__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold170 rf.registers\[12\]\[8\] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 rf.registers\[19\]\[5\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 rf.registers\[1\]\[30\] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4527__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_31_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8481__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7825__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5868__B1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7126__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6030__A _1634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4766__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4518__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5090_ rf.registers\[28\]\[17\] rf.registers\[29\]\[17\] rf.registers\[30\]\[17\]
+ rf.registers\[31\]\[17\] _1689_ _1693_ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5080__S _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5191__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6045__B1 _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7800_ net656 _3489_ _3855_ VGND VGND VPWR VPWR _3862_ sky130_fd_sc_hd__mux2_1
X_8780_ clknet_leaf_45_clk _0964_ VGND VGND VPWR VPWR rf.registers\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5992_ _2347_ _2622_ VGND VGND VPWR VPWR _2732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7731_ _3825_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__clkbuf_1
X_4943_ _1696_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7545__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7662_ net1069 _3487_ _3783_ VGND VGND VPWR VPWR _3789_ sky130_fd_sc_hd__mux2_1
X_4874_ rf.registers\[4\]\[18\] rf.registers\[5\]\[18\] rf.registers\[6\]\[18\] rf.registers\[7\]\[18\]
+ net132 _1175_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__mux4_1
XANTENNA__6205__A _1958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6613_ _3062_ net1065 _3206_ VGND VGND VPWR VPWR _3216_ sky130_fd_sc_hd__mux2_1
X_9401_ clknet_leaf_20_clk _0561_ VGND VGND VPWR VPWR rf.registers\[24\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7593_ _3752_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_119_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4454__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6544_ _3178_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__clkbuf_1
X_9332_ clknet_leaf_38_clk _0492_ VGND VGND VPWR VPWR rf.registers\[21\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9263_ clknet_leaf_10_clk _0423_ VGND VGND VPWR VPWR rf.registers\[23\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6475_ net28 VGND VGND VPWR VPWR _3139_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5859__B1 _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8214_ _4081_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__clkbuf_1
X_5426_ rf.registers\[16\]\[11\] rf.registers\[17\]\[11\] rf.registers\[18\]\[11\]
+ rf.registers\[19\]\[11\] _1675_ _1692_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__mux4_1
X_9194_ clknet_leaf_64_clk _0354_ VGND VGND VPWR VPWR rf.registers\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4757__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8145_ net216 _3493_ _4036_ VGND VGND VPWR VPWR _4045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8566__S _3006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5357_ _1702_ VGND VGND VPWR VPWR _2113_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_7_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A1_N _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4308_ _1062_ _1063_ _1035_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__mux2_1
X_8076_ _4008_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__clkbuf_1
X_5288_ _1684_ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__buf_4
X_7027_ _3436_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5182__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6814__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8978_ clknet_leaf_42_clk _0138_ VGND VGND VPWR VPWR rf.registers\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7929_ _3930_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_26_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4693__S0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7645__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5165__S _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4748__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7380__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4509__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6724__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4684__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6025__A _1874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7555__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4590_ _1344_ _1345_ _1259_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold906 rf.registers\[29\]\[2\] VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold917 rf.registers\[15\]\[3\] VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold928 rf.registers\[0\]\[3\] VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold939 rf.registers\[26\]\[25\] VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__dlygate4sd3_1
X_6260_ _2984_ _2985_ VGND VGND VPWR VPWR _2986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5211_ rf.registers\[24\]\[27\] rf.registers\[25\]\[27\] rf.registers\[26\]\[27\]
+ rf.registers\[27\]\[27\] _1767_ _1768_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__mux4_1
XANTENNA__8386__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6191_ _1996_ _2903_ _2919_ VGND VGND VPWR VPWR _2920_ sky130_fd_sc_hd__o21ba_1
XANTENNA__7290__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5142_ _1897_ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5073_ _1824_ _1825_ _1826_ _1827_ _1713_ _1828_ VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__mux4_1
XANTENNA__5164__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5104__A _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8901_ clknet_leaf_54_clk _0061_ VGND VGND VPWR VPWR rf.registers\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6634__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8832_ clknet_leaf_68_clk _1016_ VGND VGND VPWR VPWR rf.registers\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4943__A _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5975_ _2573_ _2591_ VGND VGND VPWR VPWR _2716_ sky130_fd_sc_hd__and2_1
X_8763_ clknet_leaf_21_clk _0947_ VGND VGND VPWR VPWR rf.registers\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4675__S0 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7714_ _3816_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7518__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4926_ rf.registers\[20\]\[23\] rf.registers\[21\]\[23\] rf.registers\[22\]\[23\]
+ rf.registers\[23\]\[23\] _1676_ _1681_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__mux4_1
X_8694_ clknet_leaf_24_clk _0878_ VGND VGND VPWR VPWR rf.registers\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7645_ net828 _3470_ _3772_ VGND VGND VPWR VPWR _3780_ sky130_fd_sc_hd__mux2_1
X_4857_ _1190_ _1612_ _1205_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7576_ _3743_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4788_ rf.registers\[16\]\[10\] rf.registers\[17\]\[10\] rf.registers\[18\]\[10\]
+ rf.registers\[19\]\[10\] net93 _1043_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__mux4_2
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9315_ clknet_leaf_68_clk _0475_ VGND VGND VPWR VPWR rf.registers\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6527_ net558 _3116_ _3168_ VGND VGND VPWR VPWR _3170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8494__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9246_ clknet_leaf_73_clk _0406_ VGND VGND VPWR VPWR rf.registers\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6458_ _3127_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__clkbuf_1
X_5409_ rf.registers\[20\]\[12\] rf.registers\[21\]\[12\] rf.registers\[22\]\[12\]
+ rf.registers\[23\]\[12\] _2113_ _2114_ VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__mux4_1
XANTENNA__8296__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9177_ clknet_leaf_20_clk _0337_ VGND VGND VPWR VPWR rf.registers\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6389_ _3079_ net1008 _3065_ VGND VGND VPWR VPWR _3080_ sky130_fd_sc_hd__mux2_1
X_8128_ _4024_ VGND VGND VPWR VPWR _4036_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8059_ _3999_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7757__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4666__S0 net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7375__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8060__A _3988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4969__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5091__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8485__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_53_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6454__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4975__A1_N _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5760_ _2481_ _2484_ _2480_ VGND VGND VPWR VPWR _2512_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_17_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4711_ _1465_ _1466_ _1036_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5691_ _2441_ _2444_ _2040_ VGND VGND VPWR VPWR _2445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7430_ _3666_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4642_ _1392_ _1394_ _1397_ _1078_ _1057_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7361_ _3025_ net836 _3628_ VGND VGND VPWR VPWR _3630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4573_ _1189_ _1328_ _1078_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__a21o_1
Xhold703 rf.registers\[12\]\[9\] VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd3_1
X_6312_ _3027_ net594 _3023_ VGND VGND VPWR VPWR _3028_ sky130_fd_sc_hd__mux2_1
Xhold714 rf.registers\[31\]\[2\] VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd3_1
X_9100_ clknet_leaf_46_clk _0260_ VGND VGND VPWR VPWR rf.registers\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold725 rf.registers\[27\]\[3\] VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd3_1
X_7292_ _3025_ net383 _3591_ VGND VGND VPWR VPWR _3593_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold736 rf.registers\[31\]\[10\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 rf.registers\[15\]\[6\] VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold758 rf.registers\[22\]\[3\] VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd3_1
X_9031_ clknet_leaf_66_clk _0191_ VGND VGND VPWR VPWR rf.registers\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6243_ _2420_ _2968_ _2501_ VGND VGND VPWR VPWR _2969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold769 rf.registers\[8\]\[28\] VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8228__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6174_ _1996_ _2903_ VGND VGND VPWR VPWR _2904_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_71_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5125_ _1720_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5056_ rf.registers\[8\]\[18\] rf.registers\[9\]\[18\] rf.registers\[10\]\[18\] rf.registers\[11\]\[18\]
+ _1689_ _1693_ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_127_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4896__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6364__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8815_ clknet_leaf_29_clk _0999_ VGND VGND VPWR VPWR rf.registers\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4648__S0 _1104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8746_ clknet_leaf_7_clk _0930_ VGND VGND VPWR VPWR rf.registers\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5958_ _2104_ _2696_ _2700_ VGND VGND VPWR VPWR _2701_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_80_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4909_ _1664_ _1060_ _1084_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__or3_1
X_8677_ clknet_leaf_61_clk _0861_ VGND VGND VPWR VPWR rf.registers\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5889_ _2246_ _2616_ _2634_ VGND VGND VPWR VPWR _2635_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5708__S _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4612__S _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7628_ _3770_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5073__S0 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7559_ _3087_ net888 _3699_ VGND VGND VPWR VPWR _3734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4820__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9229_ clknet_leaf_44_clk _0389_ VGND VGND VPWR VPWR rf.registers\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6539__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5376__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold63 rf.registers\[5\]\[9\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 rf.registers\[9\]\[13\] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 rf.registers\[7\]\[6\] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5453__A1 _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold96 rf.registers\[19\]\[10\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4887__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4639__S0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_119_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5845__C _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_5 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8458__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_128_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7130__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5589__A _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer17 _1315_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_109_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6930_ _3384_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer28 _2712_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer39 _1416_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_13_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6861_ net1009 _3107_ _3340_ VGND VGND VPWR VPWR _3348_ sky130_fd_sc_hd__mux2_1
X_8600_ clknet_leaf_26_clk _0784_ VGND VGND VPWR VPWR rf.registers\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5812_ _2559_ _2560_ VGND VGND VPWR VPWR _2561_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_122_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6792_ _3311_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__clkbuf_1
X_9580_ clknet_leaf_45_clk _0740_ VGND VGND VPWR VPWR rf.registers\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6944__A1 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8531_ net344 net44 _4244_ VGND VGND VPWR VPWR _4249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5743_ _2040_ _2335_ VGND VGND VPWR VPWR _2495_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5528__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4432__S _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8462_ net669 net43 _4205_ VGND VGND VPWR VPWR _4213_ sky130_fd_sc_hd__mux2_1
X_5674_ _1168_ _2230_ VGND VGND VPWR VPWR _2428_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7413_ _3077_ net1123 _3650_ VGND VGND VPWR VPWR _3657_ sky130_fd_sc_hd__mux2_1
X_4625_ rf.registers\[12\]\[24\] rf.registers\[13\]\[24\] rf.registers\[14\]\[24\]
+ rf.registers\[15\]\[24\] _1351_ _1352_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8393_ _4176_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7743__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7344_ _3077_ net1084 _3613_ VGND VGND VPWR VPWR _3620_ sky130_fd_sc_hd__mux2_1
Xhold500 rf.registers\[2\]\[22\] VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 rf.registers\[14\]\[26\] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ rf.registers\[0\]\[27\] rf.registers\[1\]\[27\] rf.registers\[2\]\[27\] rf.registers\[3\]\[27\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__mux4_1
Xhold522 rf.registers\[23\]\[7\] VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold533 rf.registers\[2\]\[25\] VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold544 rf.registers\[27\]\[28\] VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 rf.registers\[7\]\[13\] VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
X_7275_ _3583_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
Xhold566 rf.registers\[24\]\[3\] VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ rf.registers\[28\]\[20\] rf.registers\[29\]\[20\] rf.registers\[30\]\[20\]
+ rf.registers\[31\]\[20\] _1207_ _1208_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__mux4_1
XANTENNA__7121__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold577 rf.registers\[25\]\[7\] VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold588 rf.registers\[25\]\[15\] VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__dlygate4sd3_1
X_9014_ clknet_leaf_33_clk _0174_ VGND VGND VPWR VPWR rf.registers\[31\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6226_ _2951_ _2952_ VGND VGND VPWR VPWR _2953_ sky130_fd_sc_hd__or2b_1
Xhold599 rf.registers\[17\]\[0\] VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _1447_ _1384_ _2871_ _2741_ VGND VGND VPWR VPWR _2888_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5108_ rf.registers\[20\]\[16\] rf.registers\[21\]\[16\] rf.registers\[22\]\[16\]
+ rf.registers\[23\]\[16\] _1705_ _1708_ VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__mux4_1
X_6088_ _2040_ _2797_ VGND VGND VPWR VPWR _2823_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_142_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6632__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5039_ rf.registers\[0\]\[20\] rf.registers\[1\]\[20\] rf.registers\[2\]\[20\] rf.registers\[3\]\[20\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8729_ clknet_leaf_19_clk _0913_ VGND VGND VPWR VPWR rf.registers\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5173__S _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput53 net53 VGND VGND VPWR VPWR alu_out[13] sky130_fd_sc_hd__buf_2
Xoutput64 net64 VGND VGND VPWR VPWR alu_out[23] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VGND VGND VPWR VPWR alu_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5521__S1 _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7129__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7563__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4410_ _1057_ _1153_ _1157_ _1165_ _1161_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a32o_4
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5390_ rf.registers\[16\]\[13\] rf.registers\[17\]\[13\] rf.registers\[18\]\[13\]
+ rf.registers\[19\]\[13\] _1673_ _1690_ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4341_ _1095_ _1096_ _1040_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7060_ _3457_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4272_ A2[1] VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6011_ _2740_ _2730_ _2750_ _2621_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__o22a_1
XANTENNA__6907__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8394__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_145_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7962_ _3947_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5512__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5968__A2 _1480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6913_ _3155_ _3302_ VGND VGND VPWR VPWR _3375_ sky130_fd_sc_hd__nor2_4
XFILLER_0_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7893_ _3011_ net967 _3902_ VGND VGND VPWR VPWR _3911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7738__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6642__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4951__A _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6917__A1 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6844_ _3338_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9563_ clknet_leaf_21_clk _0723_ VGND VGND VPWR VPWR rf.registers\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6775_ _3301_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8514_ net728 net14 _3007_ VGND VGND VPWR VPWR _4240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5726_ _2039_ _2478_ VGND VGND VPWR VPWR _2479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9494_ clknet_leaf_33_clk _0654_ VGND VGND VPWR VPWR rf.registers\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5028__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8445_ _4203_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5657_ net1169 _2411_ _1145_ VGND VGND VPWR VPWR _2412_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7473__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4608_ _1362_ _1363_ _1190_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ _2341_ _2342_ VGND VGND VPWR VPWR _2343_ sky130_fd_sc_hd__and2b_1
X_8376_ net385 _3452_ _4132_ VGND VGND VPWR VPWR _4167_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold330 rf.registers\[16\]\[16\] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
X_7327_ _3060_ net246 _3602_ VGND VGND VPWR VPWR _3611_ sky130_fd_sc_hd__mux2_1
Xhold341 rf.registers\[28\]\[31\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ rf.registers\[12\]\[26\] rf.registers\[13\]\[26\] rf.registers\[14\]\[26\]
+ rf.registers\[15\]\[26\] net1156 _1279_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__mux4_1
Xhold352 rf.registers\[10\]\[31\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 rf.registers\[10\]\[30\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 rf.registers\[18\]\[5\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold385 rf.registers\[18\]\[21\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 rf.registers\[18\]\[6\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
X_7258_ _3574_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
X_6209_ _2875_ _2892_ VGND VGND VPWR VPWR _2937_ sky130_fd_sc_hd__nor2_1
X_7189_ net577 _3493_ _3528_ VGND VGND VPWR VPWR _3537_ sky130_fd_sc_hd__mux2_1
Xhold1030 rf.registers\[15\]\[31\] VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6605__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1041 rf.registers\[26\]\[26\] VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 rf.registers\[27\]\[4\] VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4337__S _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1063 rf.registers\[29\]\[15\] VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5503__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__5957__A _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6552__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5041__C1 _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5019__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_5_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8479__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer8 _2657_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_133_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4800__S _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5647__A1 _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output49_A net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5867__A _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4890_ _1643_ _1644_ _1645_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__mux2_1
XANTENNA__8243__A _4096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6560_ net745 _3009_ _3179_ VGND VGND VPWR VPWR _3187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_671 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5511_ rf.registers\[4\]\[6\] rf.registers\[5\]\[6\] rf.registers\[6\]\[6\] rf.registers\[7\]\[6\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2267_ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6491_ net331 _3011_ _3135_ VGND VGND VPWR VPWR _3149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5442_ rf.registers\[20\]\[10\] rf.registers\[21\]\[10\] rf.registers\[22\]\[10\]
+ rf.registers\[23\]\[10\] _2050_ _2052_ VGND VGND VPWR VPWR _2198_ sky130_fd_sc_hd__mux4_1
X_8230_ net165 _3442_ _4083_ VGND VGND VPWR VPWR _4090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5430__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5373_ rf.registers\[24\]\[14\] rf.registers\[25\]\[14\] rf.registers\[26\]\[14\]
+ rf.registers\[27\]\[14\] _1674_ _1691_ VGND VGND VPWR VPWR _2129_ sky130_fd_sc_hd__mux4_1
X_8161_ _4053_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4324_ rf.registers\[0\]\[5\] rf.registers\[1\]\[5\] rf.registers\[2\]\[5\] rf.registers\[3\]\[5\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7112_ _3492_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_8092_ net596 _3508_ _4011_ VGND VGND VPWR VPWR _4017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7043_ _3445_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4946__A _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8994_ clknet_leaf_59_clk _0154_ VGND VGND VPWR VPWR rf.registers\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7945_ net465 _3497_ _3938_ VGND VGND VPWR VPWR _3939_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7876_ _3879_ VGND VGND VPWR VPWR _3902_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6827_ net839 _3141_ _3326_ VGND VGND VPWR VPWR _3330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9546_ clknet_leaf_7_clk _0706_ VGND VGND VPWR VPWR rf.registers\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6758_ _3071_ net682 _3289_ VGND VGND VPWR VPWR _3293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5709_ _2460_ _2461_ _2252_ VGND VGND VPWR VPWR _2462_ sky130_fd_sc_hd__mux2_1
X_9477_ clknet_leaf_52_clk _0637_ VGND VGND VPWR VPWR rf.registers\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6689_ _3256_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8428_ net249 _3504_ _4191_ VGND VGND VPWR VPWR _4195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8359_ _4158_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5017__A _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold160 rf.registers\[11\]\[29\] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 rf.registers\[11\]\[25\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 rf.registers\[17\]\[14\] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 rf.registers\[7\]\[27\] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7251__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5801__B2 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4368__B2 _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4530__S _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8002__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6311__A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5412__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7841__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6457__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6293__A1 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5479__S0 _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5991_ _1111_ _2335_ VGND VGND VPWR VPWR _2731_ sky130_fd_sc_hd__nor2_2
XFILLER_0_149_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5597__A _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7730_ _3054_ net867 _3819_ VGND VGND VPWR VPWR _3825_ sky130_fd_sc_hd__mux2_1
X_4942_ _1687_ _1695_ _1697_ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7661_ _3788_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4873_ _1214_ _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__nand2_1
X_9400_ clknet_leaf_27_clk _0560_ VGND VGND VPWR VPWR rf.registers\[24\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6612_ _3215_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7592_ _3052_ net605 _3747_ VGND VGND VPWR VPWR _3752_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4454__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9331_ clknet_leaf_35_clk _0491_ VGND VGND VPWR VPWR rf.registers\[21\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6543_ net611 _3132_ _3168_ VGND VGND VPWR VPWR _3178_ sky130_fd_sc_hd__mux2_1
XANTENNA__5536__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9262_ clknet_leaf_42_clk _0422_ VGND VGND VPWR VPWR rf.registers\[23\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6474_ _3138_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8213_ net213 _3493_ _4072_ VGND VGND VPWR VPWR _4081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5425_ rf.registers\[28\]\[11\] rf.registers\[29\]\[11\] rf.registers\[30\]\[11\]
+ rf.registers\[31\]\[11\] _1675_ _1692_ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__mux4_1
X_9193_ clknet_leaf_49_clk _0353_ VGND VGND VPWR VPWR rf.registers\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7751__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5356_ _1712_ _2111_ VGND VGND VPWR VPWR _2112_ sky130_fd_sc_hd__or2_1
X_8144_ _4044_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4307_ rf.registers\[16\]\[5\] rf.registers\[17\]\[5\] rf.registers\[18\]\[5\] rf.registers\[19\]\[5\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__mux4_1
X_5287_ rf.registers\[16\]\[3\] rf.registers\[17\]\[3\] rf.registers\[18\]\[3\] rf.registers\[19\]\[3\]
+ _1674_ _1691_ VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__mux4_1
X_8075_ net224 _3491_ _4000_ VGND VGND VPWR VPWR _4008_ sky130_fd_sc_hd__mux2_1
X_7026_ net646 _3134_ _3435_ VGND VGND VPWR VPWR _3436_ sky130_fd_sc_hd__mux2_1
XANTENNA__4295__B1 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8977_ clknet_leaf_40_clk _0137_ VGND VGND VPWR VPWR rf.registers\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7198__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4593__B_N _1348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7928_ net155 _3481_ _3927_ VGND VGND VPWR VPWR _3930_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4693__S1 _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7859_ _3893_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7926__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9529_ clknet_leaf_19_clk _0689_ VGND VGND VPWR VPWR rf.registers\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6131__A _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6275__A1 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8492__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4381__S0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7775__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4684__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold907 rf.registers\[27\]\[29\] VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold918 rf.registers\[31\]\[29\] VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold929 rf.registers\[15\]\[28\] VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7571__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5210_ rf.registers\[28\]\[27\] rf.registers\[29\]\[27\] rf.registers\[30\]\[27\]
+ rf.registers\[31\]\[27\] _1767_ _1768_ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__mux4_1
X_6190_ _2875_ net136 _2892_ _2904_ _2890_ VGND VGND VPWR VPWR _2919_ sky130_fd_sc_hd__o311a_1
XFILLER_0_110_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5141_ _1693_ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__buf_4
X_5072_ _1716_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__buf_4
X_8900_ clknet_leaf_51_clk _0060_ VGND VGND VPWR VPWR rf.registers\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6915__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8831_ clknet_leaf_68_clk _1015_ VGND VGND VPWR VPWR rf.registers\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8762_ clknet_leaf_18_clk _0946_ VGND VGND VPWR VPWR rf.registers\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5974_ _2707_ _2709_ _2715_ _2621_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__o22a_2
X_7713_ _3037_ net951 _3808_ VGND VGND VPWR VPWR _3816_ sky130_fd_sc_hd__mux2_1
XANTENNA__4675__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4925_ _1680_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__clkbuf_4
X_8693_ clknet_leaf_32_clk _0877_ VGND VGND VPWR VPWR rf.registers\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6650__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5529__B1 _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7644_ _3779_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4856_ rf.registers\[0\]\[19\] rf.registers\[1\]\[19\] rf.registers\[2\]\[19\] rf.registers\[3\]\[19\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_30_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7575_ _3035_ net969 _3736_ VGND VGND VPWR VPWR _3743_ sky130_fd_sc_hd__mux2_1
X_4787_ rf.registers\[20\]\[10\] rf.registers\[21\]\[10\] rf.registers\[22\]\[10\]
+ rf.registers\[23\]\[10\] net93 _1043_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__mux4_2
XFILLER_0_90_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7047__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9314_ clknet_leaf_59_clk _0474_ VGND VGND VPWR VPWR rf.registers\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6526_ _3169_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9245_ clknet_leaf_13_clk _0405_ VGND VGND VPWR VPWR rf.registers\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6457_ net291 _3126_ _3114_ VGND VGND VPWR VPWR _3127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7481__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5408_ rf.registers\[16\]\[12\] rf.registers\[17\]\[12\] rf.registers\[18\]\[12\]
+ rf.registers\[19\]\[12\] _2113_ _2114_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9176_ clknet_leaf_12_clk _0336_ VGND VGND VPWR VPWR rf.registers\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6388_ net33 VGND VGND VPWR VPWR _3079_ sky130_fd_sc_hd__clkbuf_2
X_8127_ _4035_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__clkbuf_1
X_5339_ _2093_ _2094_ net3 VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8058_ net1033 _3474_ _3989_ VGND VGND VPWR VPWR _3999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7009_ net205 _3118_ _3424_ VGND VGND VPWR VPWR _3427_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4363__S0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6825__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4345__S _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4666__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7656__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5965__A _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6560__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5176__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5091__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8487__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5884__B_N _1542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6735__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4327__A2_N _1070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6420__A1 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ rf.registers\[16\]\[13\] rf.registers\[17\]\[13\] rf.registers\[18\]\[13\]
+ rf.registers\[19\]\[13\] net126 _1029_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6470__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5690_ _2442_ _2443_ _2252_ VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__mux2_2
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4641_ _1395_ _1396_ _1040_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7360_ _3629_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
X_4572_ rf.registers\[12\]\[31\] rf.registers\[13\]\[31\] rf.registers\[14\]\[31\]
+ rf.registers\[15\]\[31\] _1324_ _1325_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6311_ net36 VGND VGND VPWR VPWR _3027_ sky130_fd_sc_hd__clkbuf_2
Xhold704 rf.registers\[29\]\[30\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold715 rf.registers\[23\]\[21\] VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 rf.registers\[30\]\[25\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd3_1
X_7291_ _3592_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold737 rf.registers\[30\]\[11\] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9030_ clknet_leaf_0_clk _0190_ VGND VGND VPWR VPWR rf.registers\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold748 rf.registers\[4\]\[28\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 rf.registers\[14\]\[1\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd3_1
X_6242_ _2498_ _2967_ _2327_ VGND VGND VPWR VPWR _2968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6173_ net1162 _2902_ VGND VGND VPWR VPWR _2903_ sky130_fd_sc_hd__xnor2_1
X_5124_ _1804_ _1878_ _1879_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__mux2_2
X_5055_ _1807_ _1810_ _1697_ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_49_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_127_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4896__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8814_ clknet_leaf_44_clk _0998_ VGND VGND VPWR VPWR rf.registers\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6411__A1 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4648__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8745_ clknet_leaf_64_clk _0929_ VGND VGND VPWR VPWR rf.registers\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_5957_ _2104_ _2699_ VGND VGND VPWR VPWR _2700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5785__A _1059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6380__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4908_ net47 VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__inv_2
X_8676_ clknet_leaf_62_clk _0860_ VGND VGND VPWR VPWR rf.registers\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_5888_ _2229_ _2597_ _2616_ _2246_ VGND VGND VPWR VPWR _2634_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7627_ _3087_ net423 _3735_ VGND VGND VPWR VPWR _3770_ sky130_fd_sc_hd__mux2_1
X_4839_ _1593_ _1594_ _1287_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7911__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5073__S1 _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7558_ _3733_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
X_6509_ _3160_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4820__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7489_ _3085_ net522 _3663_ VGND VGND VPWR VPWR _3697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9228_ clknet_leaf_45_clk _0388_ VGND VGND VPWR VPWR rf.registers\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8100__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9159_ clknet_leaf_1_clk _0319_ VGND VGND VPWR VPWR rf.registers\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4584__S0 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5025__A _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4336__S0 _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold64 rf.registers\[11\]\[11\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5989__B1 _2729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold75 rf.registers\[16\]\[4\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 rf.registers\[9\]\[31\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6650__A1 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4887__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold97 rf.registers\[1\]\[6\] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4639__S1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5695__A _2080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7386__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6290__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_6 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8010__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output79_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4575__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer18 _1464_ VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer29 net110 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_109_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6860_ _3347_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8394__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5811_ _2286_ _2558_ VGND VGND VPWR VPWR _2560_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6791_ net821 _3105_ _3304_ VGND VGND VPWR VPWR _3311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7296__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8530_ _4248_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__clkbuf_1
X_5742_ _2105_ _2491_ _2493_ VGND VGND VPWR VPWR _2494_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8461_ _4212_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_98_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5673_ _2424_ _2425_ _2426_ VGND VGND VPWR VPWR _2427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7412_ _3656_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4624_ rf.registers\[8\]\[24\] rf.registers\[9\]\[24\] rf.registers\[10\]\[24\] rf.registers\[11\]\[24\]
+ _1351_ _1352_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__mux4_1
X_8392_ net255 _3468_ _4169_ VGND VGND VPWR VPWR _4176_ sky130_fd_sc_hd__mux2_1
XANTENNA__4707__B2 _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold501 rf.registers\[29\]\[6\] VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
X_7343_ _3619_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4949__A _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4555_ rf.registers\[4\]\[27\] rf.registers\[5\]\[27\] rf.registers\[6\]\[27\] rf.registers\[7\]\[27\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__mux4_1
Xhold512 rf.registers\[22\]\[2\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 rf.registers\[28\]\[14\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 rf.registers\[4\]\[25\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 rf.registers\[17\]\[7\] VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
X_7274_ _3075_ net1148 _3577_ VGND VGND VPWR VPWR _3583_ sky130_fd_sc_hd__mux2_1
Xhold556 rf.registers\[19\]\[4\] VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4486_ _1240_ _1241_ _1211_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__mux2_1
Xhold567 rf.registers\[20\]\[4\] VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 rf.registers\[11\]\[26\] VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__dlygate4sd3_1
X_9013_ clknet_leaf_31_clk _0173_ VGND VGND VPWR VPWR rf.registers\[31\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold589 rf.registers\[27\]\[5\] VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _1942_ _2950_ VGND VGND VPWR VPWR _2952_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_129_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7409__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6880__A1 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6156_ _2875_ _2885_ VGND VGND VPWR VPWR _2887_ sky130_fd_sc_hd__or2_1
XANTENNA__4318__S0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5107_ rf.registers\[16\]\[16\] rf.registers\[17\]\[16\] rf.registers\[18\]\[16\]
+ rf.registers\[19\]\[16\] _1705_ _1708_ VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__mux4_1
X_6087_ _2753_ _2821_ _1126_ VGND VGND VPWR VPWR _2822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5038_ rf.registers\[4\]\[20\] rf.registers\[5\]\[20\] rf.registers\[6\]\[20\] rf.registers\[7\]\[20\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_49_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6989_ _3416_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8728_ clknet_leaf_26_clk _0912_ VGND VGND VPWR VPWR rf.registers\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8137__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8659_ clknet_leaf_32_clk _0843_ VGND VGND VPWR VPWR rf.registers\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7934__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput54 net54 VGND VGND VPWR VPWR alu_out[14] sky130_fd_sc_hd__buf_6
Xoutput65 net65 VGND VGND VPWR VPWR alu_out[24] sky130_fd_sc_hd__buf_2
Xoutput76 net76 VGND VGND VPWR VPWR alu_out[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_19_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6314__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7887__A0 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4340_ rf.registers\[24\]\[3\] rf.registers\[25\]\[3\] rf.registers\[26\]\[3\] rf.registers\[27\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4548__S0 _1262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4271_ _1026_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__buf_12
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6010_ _2744_ _2749_ VGND VGND VPWR VPWR _2750_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7961_ net325 _3446_ _3938_ VGND VGND VPWR VPWR _3947_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5968__A3 _1464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6912_ _3374_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6923__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4720__S0 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7892_ _3910_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6843_ net931 _3017_ _3303_ VGND VGND VPWR VPWR _3338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5539__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6224__A _1942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9562_ clknet_leaf_18_clk _0722_ VGND VGND VPWR VPWR rf.registers\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6774_ _3087_ net1080 _3266_ VGND VGND VPWR VPWR _3301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8513_ _4239_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5725_ net84 _1145_ _1167_ _2411_ VGND VGND VPWR VPWR _2478_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9493_ clknet_leaf_35_clk _0653_ VGND VGND VPWR VPWR rf.registers\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5028__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8444_ net238 net38 _4168_ VGND VGND VPWR VPWR _4203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5656_ _2409_ VGND VGND VPWR VPWR _2411_ sky130_fd_sc_hd__buf_2
XFILLER_0_73_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4607_ rf.registers\[12\]\[25\] rf.registers\[13\]\[25\] rf.registers\[14\]\[25\]
+ rf.registers\[15\]\[25\] _1360_ _1361_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4787__S0 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8375_ _4166_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5587_ net82 _2124_ VGND VGND VPWR VPWR _2342_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold320 rf.registers\[21\]\[3\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
X_7326_ _3610_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
Xhold331 rf.registers\[4\]\[30\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4538_ rf.registers\[8\]\[26\] rf.registers\[9\]\[26\] rf.registers\[10\]\[26\] rf.registers\[11\]\[26\]
+ net1156 _1279_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__mux4_1
Xhold342 rf.registers\[6\]\[26\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold353 rf.registers\[8\]\[8\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 rf.registers\[13\]\[17\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 rf.registers\[19\]\[21\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4539__S0 net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7257_ _3058_ net777 _3566_ VGND VGND VPWR VPWR _3574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold386 rf.registers\[4\]\[16\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ rf.registers\[28\]\[28\] rf.registers\[29\]\[28\] rf.registers\[30\]\[28\]
+ rf.registers\[31\]\[28\] net127 _1222_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__mux4_1
Xhold397 rf.registers\[18\]\[3\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6853__A1 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6208_ _2893_ _2935_ VGND VGND VPWR VPWR _2936_ sky130_fd_sc_hd__nor2_1
X_7188_ _3536_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__9059__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6139_ _1512_ _2835_ net1160 _2658_ VGND VGND VPWR VPWR _2871_ sky130_fd_sc_hd__and4_1
Xhold1020 rf.registers\[27\]\[21\] VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 rf.registers\[28\]\[5\] VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 rf.registers\[25\]\[1\] VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 rf.registers\[8\]\[21\] VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 rf.registers\[28\]\[21\] VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6833__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8358__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7664__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5019__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer9 _1348_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__4778__S0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5184__S _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7839__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6743__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4702__S0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8349__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5867__B _2613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5510_ _1699_ _2265_ VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6490_ _3148_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5441_ _2195_ _2196_ _1711_ VGND VGND VPWR VPWR _2197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4769__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5430__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8160_ net962 _3508_ _4047_ VGND VGND VPWR VPWR _4053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5372_ rf.registers\[28\]\[14\] rf.registers\[29\]\[14\] rf.registers\[30\]\[14\]
+ rf.registers\[31\]\[14\] _1674_ _1691_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7111_ net462 _3491_ _3477_ VGND VGND VPWR VPWR _3492_ sky130_fd_sc_hd__mux2_1
X_4323_ rf.registers\[4\]\[5\] rf.registers\[5\]\[5\] rf.registers\[6\]\[5\] rf.registers\[7\]\[5\]
+ net103 _1044_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8091_ _4016_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5822__S _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7042_ net464 _3444_ _3435_ VGND VGND VPWR VPWR _3445_ sky130_fd_sc_hd__mux2_1
XANTENNA__5194__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5123__A _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8993_ clknet_leaf_57_clk _0153_ VGND VGND VPWR VPWR rf.registers\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7749__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4962__A _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7944_ _3915_ VGND VGND VPWR VPWR _3938_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7875_ _3901_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6826_ _3329_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_42_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9545_ clknet_leaf_6_clk _0705_ VGND VGND VPWR VPWR rf.registers\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6757_ _3292_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5708_ _2346_ _2351_ _2327_ VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__mux2_1
X_9476_ clknet_leaf_52_clk _0636_ VGND VGND VPWR VPWR rf.registers\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6688_ net802 _3139_ _3253_ VGND VGND VPWR VPWR _3256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8512__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8427_ _4194_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__clkbuf_1
X_5639_ _1168_ _1755_ VGND VGND VPWR VPWR _2394_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_150_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8358_ net316 _3502_ _4155_ VGND VGND VPWR VPWR _4158_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold150 rf.registers\[7\]\[12\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
X_7309_ _3601_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
Xhold161 rf.registers\[23\]\[4\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 rf.registers\[18\]\[31\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
X_8289_ _4121_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__clkbuf_1
Xhold183 rf.registers\[5\]\[15\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 rf.registers\[13\]\[13\] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4932__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6762__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6799__A _3303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7394__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5412__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8267__A0 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output61_A net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5549__A1_N _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7569__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5479__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6473__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5990_ _2041_ _2102_ VGND VGND VPWR VPWR _2730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4941_ _1696_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__buf_6
XFILLER_0_87_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5089__S _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7660_ net345 _3485_ _3783_ VGND VGND VPWR VPWR _3788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4872_ _1626_ _1627_ _1189_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6611_ _3060_ net633 _3206_ VGND VGND VPWR VPWR _3215_ sky130_fd_sc_hd__mux2_1
X_7591_ _3751_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9330_ clknet_leaf_37_clk _0490_ VGND VGND VPWR VPWR rf.registers\[21\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6542_ _3177_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9261_ clknet_leaf_41_clk _0421_ VGND VGND VPWR VPWR rf.registers\[23\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6473_ net420 _3137_ _3135_ VGND VGND VPWR VPWR _3138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8212_ _4080_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__clkbuf_1
X_5424_ rf.registers\[24\]\[11\] rf.registers\[25\]\[11\] rf.registers\[26\]\[11\]
+ rf.registers\[27\]\[11\] _1675_ _1692_ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_132_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9192_ clknet_leaf_46_clk _0352_ VGND VGND VPWR VPWR rf.registers\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8258__A0 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8143_ net761 _3491_ _4036_ VGND VGND VPWR VPWR _4044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6648__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5355_ rf.registers\[8\]\[15\] rf.registers\[9\]\[15\] rf.registers\[10\]\[15\] rf.registers\[11\]\[15\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__mux4_1
XANTENNA__4957__A _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6808__A1 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4306_ rf.registers\[20\]\[5\] rf.registers\[21\]\[5\] rf.registers\[22\]\[5\] rf.registers\[23\]\[5\]
+ net94 _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8074_ _4007_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__clkbuf_1
X_5286_ rf.registers\[20\]\[3\] rf.registers\[21\]\[3\] rf.registers\[22\]\[3\] rf.registers\[23\]\[3\]
+ _1674_ _1691_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__mux4_1
X_7025_ _3412_ VGND VGND VPWR VPWR _3435_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_52_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4295__A1 _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7479__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6383__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4692__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8976_ clknet_leaf_3_clk _0136_ VGND VGND VPWR VPWR rf.registers\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_7927_ _3929_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_26_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7858_ _3116_ net811 _3891_ VGND VGND VPWR VPWR _3893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6809_ _3320_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7789_ _3856_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9528_ clknet_leaf_17_clk _0688_ VGND VGND VPWR VPWR rf.registers\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9459_ clknet_leaf_34_clk _0619_ VGND VGND VPWR VPWR rf.registers\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7942__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6558__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5158__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4381__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6293__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5330__S0 _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8013__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold908 rf.registers\[31\]\[17\] VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 rf.registers\[28\]\[25\] VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5473__A1_N _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5140_ _1895_ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5071_ rf.registers\[20\]\[19\] rf.registers\[21\]\[19\] rf.registers\[22\]\[19\]
+ rf.registers\[23\]\[19\] _1676_ _1681_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8830_ clknet_leaf_0_clk _1014_ VGND VGND VPWR VPWR rf.registers\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8761_ clknet_leaf_19_clk _0945_ VGND VGND VPWR VPWR rf.registers\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5321__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5973_ net111 _2714_ VGND VGND VPWR VPWR _2715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7712_ _3815_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6931__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4924_ _1679_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8692_ clknet_leaf_30_clk _0876_ VGND VGND VPWR VPWR rf.registers\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5529__A1 _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7643_ net1122 _3468_ _3772_ VGND VGND VPWR VPWR _3779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4855_ _1211_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__or2_1
XANTENNA__5547__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4737__C1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7574_ _3742_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
X_4786_ _1533_ _1025_ _1541_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__o21ai_4
X_9313_ clknet_leaf_56_clk _0473_ VGND VGND VPWR VPWR rf.registers\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6525_ net716 _3113_ _3168_ VGND VGND VPWR VPWR _3169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9244_ clknet_leaf_16_clk _0404_ VGND VGND VPWR VPWR rf.registers\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6456_ net21 VGND VGND VPWR VPWR _3126_ sky130_fd_sc_hd__buf_2
Xclkload70 clknet_leaf_36_clk VGND VGND VPWR VPWR clkload70/Y sky130_fd_sc_hd__inv_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5407_ rf.registers\[28\]\[12\] rf.registers\[29\]\[12\] rf.registers\[30\]\[12\]
+ rf.registers\[31\]\[12\] _1703_ _1706_ VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9175_ clknet_leaf_23_clk _0335_ VGND VGND VPWR VPWR rf.registers\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6387_ _3078_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8126_ net326 _3474_ _4025_ VGND VGND VPWR VPWR _4035_ sky130_fd_sc_hd__mux2_1
X_5338_ rf.registers\[12\]\[1\] rf.registers\[13\]\[1\] rf.registers\[14\]\[1\] rf.registers\[15\]\[1\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _2094_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8057_ _3998_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__clkbuf_1
X_5269_ rf.registers\[12\]\[24\] rf.registers\[13\]\[24\] rf.registers\[14\]\[24\]
+ rf.registers\[15\]\[24\] _1881_ _1883_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__mux4_1
X_7008_ _3426_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5560__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4363__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4626__S _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6407__A _3092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7002__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5312__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8959_ clknet_leaf_74_clk _0119_ VGND VGND VPWR VPWR rf.registers\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6841__S _3303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7390__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6142__A _1384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8008__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6317__A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload6_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5303__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7847__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4640_ rf.registers\[0\]\[6\] rf.registers\[1\]\[6\] rf.registers\[2\]\[6\] rf.registers\[3\]\[6\]
+ net106 _1073_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__mux4_1
XANTENNA__6052__A _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6184__A1 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5931__A1 _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4571_ _1178_ _1326_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6310_ _3026_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold705 rf.registers\[25\]\[29\] VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd3_1
X_7290_ _3019_ net762 _3591_ VGND VGND VPWR VPWR _3592_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold716 rf.registers\[5\]\[29\] VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold727 rf.registers\[4\]\[21\] VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold738 rf.registers\[4\]\[26\] VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__dlygate4sd3_1
X_6241_ _2547_ VGND VGND VPWR VPWR _2967_ sky130_fd_sc_hd__inv_2
Xhold749 rf.registers\[2\]\[31\] VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6172_ _1447_ _2901_ _2871_ _2741_ VGND VGND VPWR VPWR _2902_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5123_ _1126_ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__clkbuf_4
X_5054_ _1808_ _1809_ _1739_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__mux2_1
XANTENNA__5542__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8813_ clknet_leaf_43_clk _0997_ VGND VGND VPWR VPWR rf.registers\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7757__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4970__A _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8744_ clknet_leaf_64_clk _0928_ VGND VGND VPWR VPWR rf.registers\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5956_ _2610_ _2698_ _2251_ VGND VGND VPWR VPWR _2699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4907_ _1148_ _1662_ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__nand2_1
X_8675_ clknet_leaf_68_clk _0859_ VGND VGND VPWR VPWR rf.registers\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5887_ _2632_ _2210_ VGND VGND VPWR VPWR _2633_ sky130_fd_sc_hd__xor2_1
XANTENNA__7058__A _3455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4838_ rf.registers\[12\]\[17\] rf.registers\[13\]\[17\] rf.registers\[14\]\[17\]
+ rf.registers\[15\]\[17\] _1191_ _1279_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__mux4_1
X_7626_ _3769_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7557_ _3085_ net1130 _3699_ VGND VGND VPWR VPWR _3733_ sky130_fd_sc_hd__mux2_1
X_4769_ rf.registers\[0\]\[8\] rf.registers\[1\]\[8\] rf.registers\[2\]\[8\] rf.registers\[3\]\[8\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6508_ net315 _3097_ _3157_ VGND VGND VPWR VPWR _3160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7488_ _3696_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7675__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6439_ net958 _3113_ _3114_ VGND VGND VPWR VPWR _3115_ sky130_fd_sc_hd__mux2_1
X_9227_ clknet_leaf_5_clk _0387_ VGND VGND VPWR VPWR rf.registers\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9158_ clknet_leaf_1_clk _0318_ VGND VGND VPWR VPWR rf.registers\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4584__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8109_ _4026_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__clkbuf_1
X_9089_ clknet_leaf_59_clk _0249_ VGND VGND VPWR VPWR rf.registers\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4336__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold65 rf.registers\[9\]\[12\] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5989__B2 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold76 rf.registers\[17\]\[17\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold87 rf.registers\[4\]\[12\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 rf.registers\[9\]\[4\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clone53_A _1181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6166__A1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6166__B2 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8498__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_7 _3022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4575__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer19 _1635_ VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_109_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7577__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5810_ _2286_ _2558_ VGND VGND VPWR VPWR _2559_ sky130_fd_sc_hd__and2_1
X_6790_ _3310_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5741_ _2250_ _2255_ _2492_ _2373_ VGND VGND VPWR VPWR _2493_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_33_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8460_ net515 net42 _4205_ VGND VGND VPWR VPWR _4212_ sky130_fd_sc_hd__mux2_1
X_5672_ _1879_ VGND VGND VPWR VPWR _2426_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_98_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7411_ _3075_ net1021 _3650_ VGND VGND VPWR VPWR _3656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4623_ _1214_ _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__nor2_1
X_8391_ _4175_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7342_ _3075_ net926 _3613_ VGND VGND VPWR VPWR _3619_ sky130_fd_sc_hd__mux2_1
XANTENNA__8201__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4554_ _1254_ _1309_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__nor2_1
Xhold502 rf.registers\[2\]\[27\] VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold513 rf.registers\[5\]\[21\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 rf.registers\[18\]\[25\] VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
X_7273_ _3582_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
Xhold535 rf.registers\[5\]\[20\] VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
X_4485_ rf.registers\[16\]\[20\] rf.registers\[17\]\[20\] rf.registers\[18\]\[20\]
+ rf.registers\[19\]\[20\] _1207_ _1208_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__mux4_1
Xhold546 rf.registers\[20\]\[26\] VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold557 rf.registers\[27\]\[10\] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5126__A _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5668__B1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9012_ clknet_leaf_42_clk _0172_ VGND VGND VPWR VPWR rf.registers\[31\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold568 rf.registers\[18\]\[26\] VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 rf.registers\[14\]\[7\] VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _1942_ _2950_ VGND VGND VPWR VPWR _2951_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6656__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6155_ _2863_ _2870_ _2886_ _2408_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__o22a_2
XANTENNA__4965__A _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5106_ rf.registers\[28\]\[16\] rf.registers\[29\]\[16\] rf.registers\[30\]\[16\]
+ rf.registers\[31\]\[16\] _1720_ _1723_ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__mux4_1
XANTENNA__8082__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4318__S1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6086_ _2790_ _2820_ _1146_ VGND VGND VPWR VPWR _2821_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ _1712_ _1792_ _1716_ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__a21o_1
XANTENNA__4643__A1 _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7487__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6988_ net375 _3097_ _3413_ VGND VGND VPWR VPWR _3416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8727_ clknet_leaf_26_clk _0911_ VGND VGND VPWR VPWR rf.registers\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5939_ _2504_ _2671_ _2682_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__a21oi_2
XFILLER_0_153_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6148__A1 _1731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8658_ clknet_leaf_25_clk _0842_ VGND VGND VPWR VPWR rf.registers\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7609_ _3069_ net1149 _3758_ VGND VGND VPWR VPWR _3761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8589_ clknet_leaf_43_clk _0773_ VGND VGND VPWR VPWR rf.registers\[22\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5872__A1_N _2229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput55 net55 VGND VGND VPWR VPWR alu_out[15] sky130_fd_sc_hd__buf_2
Xoutput66 net66 VGND VGND VPWR VPWR alu_out[25] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VGND VGND VPWR VPWR alu_out[6] sky130_fd_sc_hd__buf_4
XANTENNA__6566__S _3156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8073__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4814__S _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7584__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4493__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7426__A _3663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8021__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7639__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7860__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4270_ A2[0] VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__buf_12
XANTENNA__4548__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6476__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7811__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7960_ _3946_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6911_ net226 _3017_ _3339_ VGND VGND VPWR VPWR _3374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4720__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7891_ _3009_ net805 _3902_ VGND VGND VPWR VPWR _3910_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_59_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6842_ _3337_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6773_ _3300_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__clkbuf_1
X_9561_ clknet_leaf_18_clk _0721_ VGND VGND VPWR VPWR rf.registers\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4484__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5724_ _2468_ _2476_ VGND VGND VPWR VPWR _2477_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8512_ net1034 net38 _4204_ VGND VGND VPWR VPWR _4239_ sky130_fd_sc_hd__mux2_1
XANTENNA__7327__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9492_ clknet_leaf_38_clk _0652_ VGND VGND VPWR VPWR rf.registers\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5655_ _1145_ net1169 _2409_ VGND VGND VPWR VPWR _2410_ sky130_fd_sc_hd__or3_1
X_8443_ _4202_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4606_ rf.registers\[8\]\[25\] rf.registers\[9\]\[25\] rf.registers\[10\]\[25\] rf.registers\[11\]\[25\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8374_ net711 _3450_ _4132_ VGND VGND VPWR VPWR _4166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5586_ _1758_ _1874_ _1839_ VGND VGND VPWR VPWR _2341_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4787__S1 _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold310 rf.registers\[2\]\[2\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7325_ _3058_ net990 _3602_ VGND VGND VPWR VPWR _3610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4537_ _1198_ _1292_ _1071_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__a21o_1
Xhold321 rf.registers\[5\]\[22\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 rf.registers\[11\]\[12\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 rf.registers\[27\]\[18\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold354 rf.registers\[17\]\[2\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7256_ _3573_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
Xhold365 rf.registers\[15\]\[25\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 rf.registers\[3\]\[13\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ _1218_ _1223_ _1178_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__mux2_1
XANTENNA__4539__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold387 rf.registers\[9\]\[28\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 rf.registers\[4\]\[22\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _2904_ _2918_ VGND VGND VPWR VPWR _2935_ sky130_fd_sc_hd__nand2_1
XANTENNA__6386__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7187_ net208 _3491_ _3528_ VGND VGND VPWR VPWR _3536_ sky130_fd_sc_hd__mux2_1
X_4399_ rf.registers\[24\]\[0\] rf.registers\[25\]\[0\] rf.registers\[26\]\[0\] rf.registers\[27\]\[0\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__mux4_1
X_6138_ _2504_ _2865_ _2869_ VGND VGND VPWR VPWR _2870_ sky130_fd_sc_hd__or3_1
Xhold1010 rf.registers\[21\]\[14\] VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 rf.registers\[21\]\[0\] VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1032 rf.registers\[31\]\[24\] VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 rf.registers\[14\]\[19\] VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 rf.registers\[30\]\[5\] VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6069_ net105 _2804_ VGND VGND VPWR VPWR _2805_ sky130_fd_sc_hd__xor2_1
Xhold1065 rf.registers\[20\]\[28\] VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4475__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7945__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5041__B2 _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_86_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4778__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6296__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4702__S1 _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5375__S _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5440_ rf.registers\[28\]\[10\] rf.registers\[29\]\[10\] rf.registers\[30\]\[10\]
+ rf.registers\[31\]\[10\] _1674_ _1691_ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4769__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5371_ _2125_ _2126_ _2044_ VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7590__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7110_ net22 VGND VGND VPWR VPWR _3491_ sky130_fd_sc_hd__buf_2
X_4322_ _1050_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__clkbuf_8
X_8090_ net864 _3506_ _4011_ VGND VGND VPWR VPWR _4016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7041_ net33 VGND VGND VPWR VPWR _3444_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5194__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8992_ clknet_leaf_60_clk _0152_ VGND VGND VPWR VPWR rf.registers\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7943_ _3937_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6235__A _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7874_ _3132_ net759 _3891_ VGND VGND VPWR VPWR _3901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6825_ net590 _3139_ _3326_ VGND VGND VPWR VPWR _3329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6220__B1 _2737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9544_ clknet_leaf_65_clk _0704_ VGND VGND VPWR VPWR rf.registers\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6756_ _3069_ net1025 _3289_ VGND VGND VPWR VPWR _3292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5707_ _2402_ _2343_ _2327_ VGND VGND VPWR VPWR _2460_ sky130_fd_sc_hd__mux2_1
X_9475_ clknet_leaf_60_clk _0635_ VGND VGND VPWR VPWR rf.registers\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6687_ _3255_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5285__S _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8426_ net852 _3502_ _4191_ VGND VGND VPWR VPWR _4194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7720__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5638_ _2391_ _2392_ VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_150_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5569_ _1839_ _2324_ VGND VGND VPWR VPWR _2325_ sky130_fd_sc_hd__nand2_1
X_8357_ _4157_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold140 rf.registers\[5\]\[2\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7308_ _3041_ net1121 _3591_ VGND VGND VPWR VPWR _3601_ sky130_fd_sc_hd__mux2_1
Xhold151 rf.registers\[9\]\[9\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold162 rf.registers\[24\]\[31\] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 rf.registers\[12\]\[6\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
X_8288_ _3137_ net995 _4119_ VGND VGND VPWR VPWR _4121_ sky130_fd_sc_hd__mux2_1
Xhold184 rf.registers\[26\]\[18\] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 rf.registers\[1\]\[5\] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
X_7239_ _3564_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7005__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4932__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4696__S0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4448__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7675__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6514__A1 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5224__A _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output54_A net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6754__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6981__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6045__A3 _1634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4687__S0 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4940_ net4 VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4871_ rf.registers\[12\]\[18\] rf.registers\[13\]\[18\] rf.registers\[14\]\[18\]
+ rf.registers\[15\]\[18\] _1192_ _1195_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6610_ _3214_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__clkbuf_1
X_7590_ _3050_ net397 _3747_ VGND VGND VPWR VPWR _3751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6541_ net460 _3130_ _3168_ VGND VGND VPWR VPWR _3177_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9260_ clknet_leaf_50_clk _0420_ VGND VGND VPWR VPWR rf.registers\[23\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6472_ net27 VGND VGND VPWR VPWR _3137_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5423_ _2143_ _2177_ _2178_ VGND VGND VPWR VPWR _2179_ sky130_fd_sc_hd__mux2_1
X_8211_ net189 _3491_ _4072_ VGND VGND VPWR VPWR _4080_ sky130_fd_sc_hd__mux2_1
X_9191_ clknet_leaf_67_clk _0351_ VGND VGND VPWR VPWR rf.registers\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5713__C1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6929__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5833__S _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5354_ _2106_ _2107_ _2108_ _2109_ _1685_ _1696_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__mux4_1
X_8142_ _4043_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4305_ A2[1] VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__clkbuf_4
X_8073_ net562 _3489_ _4000_ VGND VGND VPWR VPWR _4007_ sky130_fd_sc_hd__mux2_1
X_5285_ _1880_ _2038_ _2040_ VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7024_ _3434_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4973__A _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8975_ clknet_leaf_9_clk _0135_ VGND VGND VPWR VPWR rf.registers\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4678__S0 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7926_ net508 _3479_ _3927_ VGND VGND VPWR VPWR _3929_ sky130_fd_sc_hd__mux2_1
XANTENNA__6992__A1 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7857_ _3892_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7495__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6808_ net642 _3122_ _3315_ VGND VGND VPWR VPWR _3320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7788_ net137 _3476_ _3855_ VGND VGND VPWR VPWR _3856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9527_ clknet_leaf_24_clk _0687_ VGND VGND VPWR VPWR rf.registers\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6739_ _3052_ net940 _3278_ VGND VGND VPWR VPWR _3283_ sky130_fd_sc_hd__mux2_1
XANTENNA__4850__S0 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9458_ clknet_leaf_29_clk _0618_ VGND VGND VPWR VPWR rf.registers\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8409_ net175 _3485_ _4180_ VGND VGND VPWR VPWR _4185_ sky130_fd_sc_hd__mux2_1
XANTENNA__6839__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9389_ clknet_leaf_40_clk _0549_ VGND VGND VPWR VPWR rf.registers\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5158__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5044__A _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6574__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4883__A _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5330__S1 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5094__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4841__S0 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold909 rf.registers\[23\]\[16\] VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6749__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7160__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5070_ rf.registers\[16\]\[19\] rf.registers\[17\]\[19\] rf.registers\[18\]\[19\]
+ rf.registers\[19\]\[19\] _1676_ _1681_ VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8760_ clknet_leaf_17_clk _0944_ VGND VGND VPWR VPWR rf.registers\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5321__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5972_ _2669_ _2689_ _2713_ VGND VGND VPWR VPWR _2714_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7711_ _3035_ net849 _3808_ VGND VGND VPWR VPWR _3815_ sky130_fd_sc_hd__mux2_1
X_4923_ _1678_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__buf_4
X_8691_ clknet_leaf_33_clk _0875_ VGND VGND VPWR VPWR rf.registers\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7642_ _3778_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_1
X_4854_ rf.registers\[4\]\[19\] rf.registers\[5\]\[19\] rf.registers\[6\]\[19\] rf.registers\[7\]\[19\]
+ net132 _1175_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7573_ _3033_ net1113 _3736_ VGND VGND VPWR VPWR _3742_ sky130_fd_sc_hd__mux2_1
X_4785_ _1537_ _1535_ _1540_ _1088_ net8 VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4832__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9312_ clknet_leaf_69_clk _0472_ VGND VGND VPWR VPWR rf.registers\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6524_ _3156_ VGND VGND VPWR VPWR _3168_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__8479__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9243_ clknet_leaf_22_clk _0403_ VGND VGND VPWR VPWR rf.registers\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6455_ _3125_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload60 clknet_leaf_39_clk VGND VGND VPWR VPWR clkload60/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload71 clknet_leaf_37_clk VGND VGND VPWR VPWR clkload71/Y sky130_fd_sc_hd__inv_6
X_5406_ rf.registers\[24\]\[12\] rf.registers\[25\]\[12\] rf.registers\[26\]\[12\]
+ rf.registers\[27\]\[12\] _2113_ _2114_ VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6386_ _3077_ net574 _3065_ VGND VGND VPWR VPWR _3078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9174_ clknet_leaf_24_clk _0334_ VGND VGND VPWR VPWR rf.registers\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5337_ rf.registers\[8\]\[1\] rf.registers\[9\]\[1\] rf.registers\[10\]\[1\] rf.registers\[11\]\[1\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__mux4_1
X_8125_ _4034_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__clkbuf_1
X_8056_ net838 _3472_ _3989_ VGND VGND VPWR VPWR _3998_ sky130_fd_sc_hd__mux2_1
X_5268_ _2020_ _2023_ _1766_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__mux2_1
X_7007_ net667 _3116_ _3424_ VGND VGND VPWR VPWR _3426_ sky130_fd_sc_hd__mux2_1
XANTENNA__8175__A _4060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5199_ rf.registers\[12\]\[28\] rf.registers\[13\]\[28\] rf.registers\[14\]\[28\]
+ rf.registers\[15\]\[28\] _1896_ _1898_ VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_145_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5560__S1 _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8403__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8958_ clknet_leaf_74_clk _0118_ VGND VGND VPWR VPWR rf.registers\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5312__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7909_ net479 _3462_ _3916_ VGND VGND VPWR VPWR _3920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8889_ clknet_leaf_20_clk _0049_ VGND VGND VPWR VPWR rf.registers\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8114__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout2_A _1172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7953__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4823__S0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7142__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5303__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5648__S _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4570_ rf.registers\[8\]\[31\] rf.registers\[9\]\[31\] rf.registers\[10\]\[31\] rf.registers\[11\]\[31\]
+ _1324_ _1325_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6479__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold706 rf.registers\[16\]\[11\] VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold717 rf.registers\[2\]\[21\] VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 rf.registers\[9\]\[15\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6240_ _2442_ _2942_ VGND VGND VPWR VPWR _2966_ sky130_fd_sc_hd__or2_1
Xhold739 rf.registers\[6\]\[6\] VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6171_ _1385_ VGND VGND VPWR VPWR _2901_ sky130_fd_sc_hd__inv_2
X_5122_ _1841_ _1876_ _1877_ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5053_ rf.registers\[24\]\[18\] rf.registers\[25\]\[18\] rf.registers\[26\]\[18\]
+ rf.registers\[27\]\[18\] _1734_ _1735_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__mux4_1
XANTENNA__5542__S1 _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8812_ clknet_leaf_46_clk _0996_ VGND VGND VPWR VPWR rf.registers\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6942__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8743_ clknet_leaf_66_clk _0927_ VGND VGND VPWR VPWR rf.registers\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5955_ _2649_ _2697_ _1803_ VGND VGND VPWR VPWR _2698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5558__S net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4906_ _1169_ _1661_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__and2_1
X_8674_ clknet_leaf_60_clk _0858_ VGND VGND VPWR VPWR rf.registers\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5886_ _1558_ _2631_ VGND VGND VPWR VPWR _2632_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7625_ _3085_ net718 _3735_ VGND VGND VPWR VPWR _3769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4837_ rf.registers\[8\]\[17\] rf.registers\[9\]\[17\] rf.registers\[10\]\[17\] rf.registers\[11\]\[17\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__mux4_1
XANTENNA__7773__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4805__S0 _1072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5383__B1 _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7556_ _3732_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4768_ rf.registers\[4\]\[8\] rf.registers\[5\]\[8\] rf.registers\[6\]\[8\] rf.registers\[7\]\[8\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6389__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6507_ _3159_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7124__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5293__S _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4699_ _1451_ _1454_ _1071_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__mux2_1
X_7487_ _3083_ net787 _3686_ VGND VGND VPWR VPWR _3696_ sky130_fd_sc_hd__mux2_1
X_9226_ clknet_leaf_7_clk _0386_ VGND VGND VPWR VPWR rf.registers\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6438_ _3092_ VGND VGND VPWR VPWR _3114_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9157_ clknet_leaf_54_clk _0317_ VGND VGND VPWR VPWR rf.registers\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6369_ _3066_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8108_ net850 _3454_ _4025_ VGND VGND VPWR VPWR _4026_ sky130_fd_sc_hd__mux2_1
X_9088_ clknet_leaf_60_clk _0248_ VGND VGND VPWR VPWR rf.registers\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8039_ _3988_ VGND VGND VPWR VPWR _3989_ sky130_fd_sc_hd__clkbuf_8
Xhold55 rf.registers\[9\]\[10\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7013__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold66 rf.registers\[1\]\[31\] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 rf.registers\[17\]\[31\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 rf.registers\[9\]\[18\] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold99 rf.registers\[8\]\[13\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6938__A1 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clone46_A _1219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5610__A1 _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5049__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7683__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6299__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4401__A _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6626__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8019__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7858__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6762__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8543__A _3006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6929__A1 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5378__S _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5740_ _2336_ _2328_ VGND VGND VPWR VPWR _2492_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_106_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5671_ _2177_ _2213_ _2363_ VGND VGND VPWR VPWR _2425_ sky130_fd_sc_hd__mux2_1
XANTENNA__6157__A2 _1384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7410_ _3655_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__clkbuf_1
X_4622_ _1376_ _1377_ _1199_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__mux2_1
X_8390_ net269 _3466_ _4169_ VGND VGND VPWR VPWR _4175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7341_ _3618_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4553_ _1307_ _1308_ _1199_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold503 rf.registers\[10\]\[12\] VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold514 rf.registers\[20\]\[25\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold525 rf.registers\[15\]\[9\] VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5117__B1 _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7272_ _3073_ rf.registers\[29\]\[24\] _3577_ VGND VGND VPWR VPWR _3582_ sky130_fd_sc_hd__mux2_1
X_4484_ rf.registers\[20\]\[20\] rf.registers\[21\]\[20\] rf.registers\[22\]\[20\]
+ rf.registers\[23\]\[20\] _1207_ _1208_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__mux4_1
Xhold536 rf.registers\[2\]\[28\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 rf.registers\[8\]\[4\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold558 rf.registers\[25\]\[28\] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
X_9011_ clknet_leaf_34_clk _0171_ VGND VGND VPWR VPWR rf.registers\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6223_ net130 _2949_ VGND VGND VPWR VPWR _2950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold569 rf.registers\[21\]\[24\] VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_115_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6154_ _2884_ _2885_ VGND VGND VPWR VPWR _2886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5105_ rf.registers\[24\]\[16\] rf.registers\[25\]\[16\] rf.registers\[26\]\[16\]
+ rf.registers\[27\]\[16\] _1705_ _1708_ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__mux4_1
X_6085_ _2398_ _2395_ VGND VGND VPWR VPWR _2820_ sky130_fd_sc_hd__nor2_1
XANTENNA__5142__A _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5036_ rf.registers\[12\]\[20\] rf.registers\[13\]\[20\] rf.registers\[14\]\[20\]
+ rf.registers\[15\]\[20\] _1719_ _1722_ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_142_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6987_ _3415_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8726_ clknet_leaf_32_clk _0910_ VGND VGND VPWR VPWR rf.registers\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5938_ _1087_ _2678_ _2681_ VGND VGND VPWR VPWR _2682_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_62_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8657_ clknet_leaf_42_clk _0841_ VGND VGND VPWR VPWR rf.registers\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5869_ net116 _2615_ VGND VGND VPWR VPWR _2616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7608_ _3760_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8588_ clknet_leaf_50_clk _0772_ VGND VGND VPWR VPWR rf.registers\[22\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5451__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7539_ _3067_ net1102 _3722_ VGND VGND VPWR VPWR _3724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5317__A _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9209_ clknet_leaf_19_clk _0369_ VGND VGND VPWR VPWR rf.registers\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6847__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput56 net56 VGND VGND VPWR VPWR alu_out[16] sky130_fd_sc_hd__buf_4
Xoutput67 net67 VGND VGND VPWR VPWR alu_out[26] sky130_fd_sc_hd__buf_2
Xoutput78 net78 VGND VGND VPWR VPWR alu_out[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_73_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4367__S _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6084__B2 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6582__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4493__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8302__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5347__B1 _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5442__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7272__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7588__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5822__A1 _2469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6910_ _3373_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__clkbuf_1
X_7890_ _3909_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__clkbuf_1
X_6841_ net963 _3015_ _3303_ VGND VGND VPWR VPWR _3337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5586__B1 _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9560_ clknet_leaf_26_clk _0720_ VGND VGND VPWR VPWR rf.registers\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6772_ _3085_ net921 _3266_ VGND VGND VPWR VPWR _3300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8511_ _4238_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4484__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5723_ _2471_ _2475_ _2040_ VGND VGND VPWR VPWR _2476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9491_ clknet_leaf_36_clk _0651_ VGND VGND VPWR VPWR rf.registers\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8442_ net336 net37 _4168_ VGND VGND VPWR VPWR _4202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5654_ _1664_ net48 VGND VGND VPWR VPWR _2409_ sky130_fd_sc_hd__nor2_1
XANTENNA__5889__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5433__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4605_ _1352_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8373_ _4165_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5585_ _2178_ _2339_ VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold300 rf.registers\[31\]\[31\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_135_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7324_ _3609_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
Xhold311 rf.registers\[19\]\[30\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_135_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4536_ rf.registers\[0\]\[26\] rf.registers\[1\]\[26\] rf.registers\[2\]\[26\] rf.registers\[3\]\[26\]
+ _1291_ _1194_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold322 rf.registers\[13\]\[25\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold333 rf.registers\[17\]\[13\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 rf.registers\[29\]\[11\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 rf.registers\[13\]\[5\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 rf.registers\[18\]\[10\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6667__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7255_ _3056_ net1024 _3566_ VGND VGND VPWR VPWR _3573_ sky130_fd_sc_hd__mux2_1
XANTENNA__4976__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4467_ rf.registers\[16\]\[28\] rf.registers\[17\]\[28\] rf.registers\[18\]\[28\]
+ rf.registers\[19\]\[28\] _1220_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__mux4_1
Xhold377 rf.registers\[25\]\[31\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold388 rf.registers\[28\]\[0\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 rf.registers\[23\]\[6\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _2932_ _2933_ VGND VGND VPWR VPWR _2934_ sky130_fd_sc_hd__nor2_1
X_4398_ rf.registers\[28\]\[0\] rf.registers\[29\]\[0\] rf.registers\[30\]\[0\] rf.registers\[31\]\[0\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__mux4_1
X_7186_ _3535_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_6137_ _2104_ _2736_ _2868_ _1086_ VGND VGND VPWR VPWR _2869_ sky130_fd_sc_hd__o211a_1
Xhold1000 rf.registers\[18\]\[23\] VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1011 rf.registers\[23\]\[25\] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 rf.registers\[27\]\[26\] VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 rf.registers\[15\]\[15\] VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 rf.registers\[22\]\[29\] VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__dlygate4sd3_1
X_6068_ _1512_ _1635_ _2658_ _2536_ VGND VGND VPWR VPWR _2804_ sky130_fd_sc_hd__a31o_1
Xhold1055 rf.registers\[10\]\[24\] VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 rf.registers\[29\]\[25\] VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__dlygate4sd3_1
X_5019_ rf.registers\[0\]\[21\] rf.registers\[1\]\[21\] rf.registers\[2\]\[21\] rf.registers\[3\]\[21\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4475__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8709_ clknet_leaf_62_clk _0893_ VGND VGND VPWR VPWR rf.registers\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8122__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4650__S _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6431__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5424__S0 _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7961__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5047__A _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5481__S _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_43_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5804__B2 _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4825__S _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5510__A _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5415__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5370_ rf.registers\[16\]\[14\] rf.registers\[17\]\[14\] rf.registers\[18\]\[14\]
+ rf.registers\[19\]\[14\] _1674_ _1691_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4321_ _1071_ _1076_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__nand2_1
XANTENNA__6487__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5391__S _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7172__A _3516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7040_ _3443_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7245__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8991_ clknet_leaf_74_clk _0151_ VGND VGND VPWR VPWR rf.registers\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7796__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__8207__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7942_ net365 _3495_ _3927_ VGND VGND VPWR VPWR _3937_ sky130_fd_sc_hd__mux2_1
XANTENNA__7111__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7873_ _3900_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6950__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6824_ _3328_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6220__A1 _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9543_ clknet_leaf_5_clk _0703_ VGND VGND VPWR VPWR rf.registers\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6755_ _3291_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5706_ _1128_ _2458_ _2421_ VGND VGND VPWR VPWR _2459_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_154_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9474_ clknet_leaf_55_clk _0634_ VGND VGND VPWR VPWR rf.registers\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_30_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
X_6686_ net1135 _3137_ _3253_ VGND VGND VPWR VPWR _3255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5406__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8425_ _4193_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__clkbuf_1
X_5637_ _1799_ _1732_ VGND VGND VPWR VPWR _2392_ sky130_fd_sc_hd__and2_1
XANTENNA__7781__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8356_ net775 _3500_ _4155_ VGND VGND VPWR VPWR _4157_ sky130_fd_sc_hd__mux2_1
X_5568_ _1842_ _2323_ VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__nor2_1
Xhold130 rf.registers\[11\]\[8\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
X_7307_ _3600_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold141 rf.registers\[4\]\[18\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4519_ _1273_ _1274_ _1211_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__mux2_1
Xhold152 rf.registers\[6\]\[9\] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
X_8287_ _4120_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7082__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5499_ _2254_ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__buf_2
Xhold163 rf.registers\[8\]\[29\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 rf.registers\[18\]\[17\] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 rf.registers\[11\]\[5\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
X_7238_ _3039_ net908 _3555_ VGND VGND VPWR VPWR _3564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold196 rf.registers\[8\]\[11\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
X_7169_ _3526_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6039__A1 _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7021__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4696__S1 _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4448__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6161__A _2015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_40_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7691__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5722__A0 _2472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4384__S0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8027__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6336__A _3022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4687__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4461__B1 _1216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7866__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6770__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4870_ rf.registers\[8\]\[18\] rf.registers\[9\]\[18\] rf.registers\[10\]\[18\] rf.registers\[11\]\[18\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6540_ _3176_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6071__A _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6471_ _3136_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8210_ _4079_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__clkbuf_1
X_5422_ _1877_ VGND VGND VPWR VPWR _2178_ sky130_fd_sc_hd__clkbuf_4
X_9190_ clknet_leaf_0_clk _0350_ VGND VGND VPWR VPWR rf.registers\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8141_ net695 _3489_ _4036_ VGND VGND VPWR VPWR _4043_ sky130_fd_sc_hd__mux2_1
X_5353_ rf.registers\[24\]\[15\] rf.registers\[25\]\[15\] rf.registers\[26\]\[15\]
+ rf.registers\[27\]\[15\] _1782_ _1680_ VGND VGND VPWR VPWR _2109_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7466__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4304_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__buf_4
X_8072_ _4006_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__clkbuf_1
X_5284_ net81 VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__clkbuf_4
X_7023_ net919 _3132_ _3424_ VGND VGND VPWR VPWR _3434_ sky130_fd_sc_hd__mux2_1
XANTENNA__7630__A _3771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8974_ clknet_leaf_43_clk _0134_ VGND VGND VPWR VPWR rf.registers\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4678__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7925_ _3928_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7856_ _3113_ net720 _3891_ VGND VGND VPWR VPWR _3892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8194__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6807_ _3319_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7787_ _3843_ VGND VGND VPWR VPWR _3855_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4999_ _1639_ _1754_ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9526_ clknet_leaf_32_clk _0686_ VGND VGND VPWR VPWR rf.registers\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6738_ _3282_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4850__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9457_ clknet_leaf_29_clk _0617_ VGND VGND VPWR VPWR rf.registers\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6669_ net181 _3120_ _3242_ VGND VGND VPWR VPWR _3246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8408_ _4184_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9388_ clknet_leaf_49_clk _0548_ VGND VGND VPWR VPWR rf.registers\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8339_ net327 _3483_ _4144_ VGND VGND VPWR VPWR _4148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5325__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6855__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4366__S0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4375__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5148__A1_N _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6590__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7932__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5094__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4841__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5934__S _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7448__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4357__S0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6671__A1 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__6423__A1 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5971_ net1166 _2688_ _2687_ VGND VGND VPWR VPWR _2713_ sky130_fd_sc_hd__o21ba_1
XANTENNA__7596__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7710_ _3814_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4922_ _1677_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__buf_4
X_8690_ clknet_leaf_27_clk _0874_ VGND VGND VPWR VPWR rf.registers\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7641_ net296 _3466_ _3772_ VGND VGND VPWR VPWR _3778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4853_ _1605_ _1608_ _1187_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7572_ _3741_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4737__B2 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4784_ _1538_ _1539_ _1107_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__mux2_1
X_9311_ clknet_leaf_73_clk _0471_ VGND VGND VPWR VPWR rf.registers\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6523_ _3167_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4832__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8220__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9242_ clknet_leaf_18_clk _0402_ VGND VGND VPWR VPWR rf.registers\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6454_ net190 _3124_ _3114_ VGND VGND VPWR VPWR _3125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload50 clknet_leaf_28_clk VGND VGND VPWR VPWR clkload50/Y sky130_fd_sc_hd__inv_8
X_5405_ _2144_ _2160_ _1800_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__a21oi_1
Xclkload61 clknet_leaf_40_clk VGND VGND VPWR VPWR clkload61/Y sky130_fd_sc_hd__clkinv_8
Xclkload72 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload72/Y sky130_fd_sc_hd__inv_12
X_9173_ clknet_leaf_32_clk _0333_ VGND VGND VPWR VPWR rf.registers\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6385_ net32 VGND VGND VPWR VPWR _3077_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5145__A _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8124_ net350 _3472_ _4025_ VGND VGND VPWR VPWR _4034_ sky130_fd_sc_hd__mux2_1
X_5336_ net3 _2091_ _1655_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__o21a_1
XANTENNA__8100__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8055_ _3997_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6675__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5267_ _2021_ _2022_ _1745_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__mux2_1
X_7006_ _3425_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
X_5198_ rf.registers\[8\]\[28\] rf.registers\[9\]\[28\] rf.registers\[10\]\[28\] rf.registers\[11\]\[28\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_145_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4673__B1 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8957_ clknet_leaf_16_clk _0117_ VGND VGND VPWR VPWR rf.registers\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7908_ _3919_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__clkbuf_1
X_8888_ clknet_leaf_27_clk _0048_ VGND VGND VPWR VPWR rf.registers\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7839_ _3097_ net672 _3880_ VGND VGND VPWR VPWR _3883_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload0 clknet_3_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4823__S1 _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9509_ clknet_leaf_61_clk _0669_ VGND VGND VPWR VPWR rf.registers\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4339__S0 _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6102__B1 _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7602__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8040__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8330__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold707 rf.registers\[29\]\[14\] VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 rf.registers\[17\]\[1\] VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold729 rf.registers\[23\]\[11\] VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6170_ _2621_ _2894_ _2900_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__o21a_1
XFILLER_0_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5121_ _1145_ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6495__S _3092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7841__A0 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6644__A1 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5052_ rf.registers\[28\]\[18\] rf.registers\[29\]\[18\] rf.registers\[30\]\[18\]
+ rf.registers\[31\]\[18\] _1734_ _1735_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8811_ clknet_leaf_4_clk _0995_ VGND VGND VPWR VPWR rf.registers\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8742_ clknet_leaf_1_clk _0926_ VGND VGND VPWR VPWR rf.registers\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8215__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6524__A _3156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5954_ _2345_ _2349_ VGND VGND VPWR VPWR _2697_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4502__S0 _1220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4905_ _1639_ _1660_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__nor2_1
X_8673_ clknet_leaf_60_clk _0857_ VGND VGND VPWR VPWR rf.registers\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5885_ _2630_ _2594_ _2593_ net121 _2595_ VGND VGND VPWR VPWR _2631_ sky130_fd_sc_hd__o41a_1
XFILLER_0_118_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7624_ _3768_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4836_ _1588_ _1589_ _1590_ _1591_ _1287_ _1078_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4805__S1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5383__A1 _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7555_ _3083_ net989 _3722_ VGND VGND VPWR VPWR _3732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4767_ _1047_ _1522_ _1037_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__o21a_1
XANTENNA__4979__A _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6506_ net330 _3095_ _3157_ VGND VGND VPWR VPWR _3159_ sky130_fd_sc_hd__mux2_1
XANTENNA__4591__C1 _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7486_ _3695_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4698_ _1452_ _1453_ _1036_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__mux2_1
X_9225_ clknet_leaf_6_clk _0385_ VGND VGND VPWR VPWR rf.registers\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6437_ net15 VGND VGND VPWR VPWR _3113_ sky130_fd_sc_hd__buf_2
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9156_ clknet_leaf_51_clk _0316_ VGND VGND VPWR VPWR rf.registers\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6368_ _3064_ net483 _3065_ VGND VGND VPWR VPWR _3066_ sky130_fd_sc_hd__mux2_1
X_8107_ _4024_ VGND VGND VPWR VPWR _4025_ sky130_fd_sc_hd__clkbuf_8
X_5319_ net3 _2074_ _1655_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__a21o_1
X_9087_ clknet_leaf_74_clk _0247_ VGND VGND VPWR VPWR rf.registers\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6299_ net434 _3017_ _3007_ VGND VGND VPWR VPWR _3018_ sky130_fd_sc_hd__mux2_1
XANTENNA__5603__A _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8038_ _3987_ _3155_ VGND VGND VPWR VPWR _3988_ sky130_fd_sc_hd__nor2_4
Xhold56 rf.registers\[9\]\[11\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 rf.registers\[0\]\[13\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 rf.registers\[24\]\[23\] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4741__S0 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold89 rf.registers\[25\]\[13\] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8388__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9331__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4653__S _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6434__A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5049__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8560__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4889__A net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5484__S _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_9 _4096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6874__A1 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4980__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7204__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4732__S0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8579__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4563__S _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8035__S _3951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8000__A0 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7874__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5670_ _2423_ _2143_ _1147_ VGND VGND VPWR VPWR _2424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4621_ rf.registers\[0\]\[24\] rf.registers\[1\]\[24\] rf.registers\[2\]\[24\] rf.registers\[3\]\[24\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__mux4_1
XANTENNA__4799__S0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5394__S _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7340_ _3073_ net1114 _3613_ VGND VGND VPWR VPWR _3618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4552_ rf.registers\[8\]\[27\] rf.registers\[9\]\[27\] rf.registers\[10\]\[27\] rf.registers\[11\]\[27\]
+ _1267_ _1268_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold504 rf.registers\[16\]\[28\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 rf.registers\[4\]\[1\] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5117__A1 _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7271_ _3581_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold526 rf.registers\[10\]\[17\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ _1215_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__buf_4
Xhold537 rf.registers\[12\]\[4\] VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold548 rf.registers\[29\]\[26\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd3_1
X_9010_ clknet_leaf_42_clk _0170_ VGND VGND VPWR VPWR rf.registers\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6865__A1 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold559 rf.registers\[6\]\[12\] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ net97 _2741_ _2930_ VGND VGND VPWR VPWR _2949_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6153_ _2879_ _2883_ _2877_ VGND VGND VPWR VPWR _2885_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6108__A_N _1779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7114__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5104_ _1168_ _1859_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6084_ _2795_ _2798_ _2803_ _2819_ _2408_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__o32a_1
X_5035_ _1686_ _1790_ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_142_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6986_ net1002 _3095_ _3413_ VGND VGND VPWR VPWR _3415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5937_ _2491_ _2591_ _2680_ VGND VGND VPWR VPWR _2681_ sky130_fd_sc_hd__a21bo_1
X_8725_ clknet_leaf_31_clk _0909_ VGND VGND VPWR VPWR rf.registers\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8656_ clknet_leaf_10_clk _0840_ VGND VGND VPWR VPWR rf.registers\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_5868_ net115 net121 _2593_ _2594_ _2595_ VGND VGND VPWR VPWR _2615_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_11_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7607_ _3067_ net1146 _3758_ VGND VGND VPWR VPWR _3760_ sky130_fd_sc_hd__mux2_1
X_4819_ rf.registers\[28\]\[16\] rf.registers\[29\]\[16\] rf.registers\[30\]\[16\]
+ rf.registers\[31\]\[16\] _1291_ _1174_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8587_ clknet_leaf_2_clk _0771_ VGND VGND VPWR VPWR rf.registers\[22\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5799_ _2546_ _2548_ _2501_ VGND VGND VPWR VPWR _2549_ sky130_fd_sc_hd__mux2_1
XANTENNA__7085__A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5451__S1 _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7538_ _3723_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7469_ _3064_ net865 _3686_ VGND VGND VPWR VPWR _3687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9208_ clknet_leaf_11_clk _0368_ VGND VGND VPWR VPWR rf.registers\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xoutput57 net57 VGND VGND VPWR VPWR alu_out[17] sky130_fd_sc_hd__buf_2
X_9139_ clknet_leaf_35_clk _0299_ VGND VGND VPWR VPWR rf.registers\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xoutput68 net68 VGND VGND VPWR VPWR alu_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput79 net79 VGND VGND VPWR VPWR alu_out[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_73_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7959__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6863__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8533__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5347__A1 _1127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5442__S1 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4412__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output77_A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6339__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4953__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4705__S0 net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6840_ _3336_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5130__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6771_ _3299_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8510_ net602 net37 _4204_ VGND VGND VPWR VPWR _4238_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5722_ _2472_ _2474_ _2251_ VGND VGND VPWR VPWR _2475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9490_ clknet_leaf_39_clk _0650_ VGND VGND VPWR VPWR rf.registers\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8441_ _4201_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__clkbuf_1
X_5653_ _2333_ VGND VGND VPWR VPWR _2408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5433__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4604_ _1351_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__buf_4
XANTENNA__4322__A _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8372_ net902 _3448_ _4155_ VGND VGND VPWR VPWR _4165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5584_ _1799_ _2098_ _2338_ VGND VGND VPWR VPWR _2339_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8288__A0 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7323_ _3056_ net1076 _3602_ VGND VGND VPWR VPWR _3609_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold301 rf.registers\[31\]\[1\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4535_ _1290_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__6948__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold312 rf.registers\[7\]\[15\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 rf.registers\[16\]\[1\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold334 rf.registers\[18\]\[7\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7254_ _3572_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
Xhold345 rf.registers\[3\]\[16\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold356 rf.registers\[19\]\[18\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
X_4466_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__buf_4
Xhold367 rf.registers\[10\]\[5\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4976__B _1731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold378 rf.registers\[0\]\[18\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 rf.registers\[20\]\[22\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
X_6205_ _1958_ _2931_ VGND VGND VPWR VPWR _2933_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4468__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7185_ net295 _3489_ _3528_ VGND VGND VPWR VPWR _3535_ sky130_fd_sc_hd__mux2_1
XANTENNA__6249__A _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4397_ _1088_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6136_ _2254_ _2801_ _2867_ _2336_ VGND VGND VPWR VPWR _2868_ sky130_fd_sc_hd__o22a_1
Xhold1001 rf.registers\[30\]\[30\] VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7779__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1012 rf.registers\[22\]\[16\] VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1023 rf.registers\[26\]\[6\] VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ _2799_ _2731_ _2802_ _2496_ VGND VGND VPWR VPWR _2803_ sky130_fd_sc_hd__a22o_1
Xhold1034 rf.registers\[21\]\[19\] VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4992__A _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1045 rf.registers\[15\]\[30\] VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 rf.registers\[29\]\[21\] VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 rf.registers\[28\]\[22\] VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__dlygate4sd3_1
X_5018_ rf.registers\[4\]\[21\] rf.registers\[5\]\[21\] rf.registers\[6\]\[21\] rf.registers\[7\]\[21\]
+ _1705_ _1708_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6969_ net820 _3002_ _3398_ VGND VGND VPWR VPWR _3405_ sky130_fd_sc_hd__mux2_1
XANTENNA__7808__A _3843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4931__S _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4785__C1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8708_ clknet_leaf_62_clk _0892_ VGND VGND VPWR VPWR rf.registers\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8403__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8639_ clknet_leaf_70_clk _0823_ VGND VGND VPWR VPWR rf.registers\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7019__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5424__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4378__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6159__A _2015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold890 rf.registers\[25\]\[17\] VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5998__A _1127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7689__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_143_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5415__S1 _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6768__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4320_ _1074_ _1075_ _1048_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4926__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8990_ clknet_leaf_74_clk _0150_ VGND VGND VPWR VPWR rf.registers\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_7941_ _3936_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5351__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4317__A _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7872_ _3130_ net746 _3891_ VGND VGND VPWR VPWR _3900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6823_ net896 _3137_ _3326_ VGND VGND VPWR VPWR _3328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9542_ clknet_leaf_5_clk _0702_ VGND VGND VPWR VPWR rf.registers\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6754_ _3067_ net1140 _3289_ VGND VGND VPWR VPWR _3291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5705_ _2455_ _2457_ _1146_ VGND VGND VPWR VPWR _2458_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_137_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9473_ clknet_leaf_56_clk _0633_ VGND VGND VPWR VPWR rf.registers\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6685_ _3254_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5406__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5636_ net82 _2034_ VGND VGND VPWR VPWR _2391_ sky130_fd_sc_hd__and2_1
X_8424_ net668 _3500_ _4191_ VGND VGND VPWR VPWR _4193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8355_ _4156_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5567_ _1728_ _2314_ _2318_ _2322_ VGND VGND VPWR VPWR _2323_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7306_ _3039_ net795 _3591_ VGND VGND VPWR VPWR _3600_ sky130_fd_sc_hd__mux2_1
Xhold120 rf.registers\[5\]\[13\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 rf.registers\[1\]\[18\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ rf.registers\[0\]\[21\] rf.registers\[1\]\[21\] rf.registers\[2\]\[21\] rf.registers\[3\]\[21\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_57_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold142 rf.registers\[20\]\[17\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
X_8286_ _3134_ net960 _4119_ VGND VGND VPWR VPWR _4120_ sky130_fd_sc_hd__mux2_1
Xhold153 rf.registers\[6\]\[1\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ net81 _1126_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__or2_2
Xhold164 rf.registers\[31\]\[18\] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
X_7237_ _3563_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
Xhold175 rf.registers\[5\]\[6\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _1078_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__clkbuf_8
Xhold186 rf.registers\[11\]\[20\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 rf.registers\[13\]\[8\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
X_7168_ net323 _3472_ _3517_ VGND VGND VPWR VPWR _3526_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _1446_ _2741_ _2836_ VGND VGND VPWR VPWR _2852_ sky130_fd_sc_hd__o21ai_1
X_7099_ net458 _3483_ _3477_ VGND VGND VPWR VPWR _3484_ sky130_fd_sc_hd__mux2_1
XANTENNA__7302__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6747__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8133__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clone21_A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6588__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4384__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8308__S _4096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7212__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5238__B1 _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5333__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4461__A1 _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_151_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6470_ net440 _3134_ _3135_ VGND VGND VPWR VPWR _3136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5421_ _2161_ _2176_ VGND VGND VPWR VPWR _2177_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5713__A1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8140_ _4042_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5352_ rf.registers\[28\]\[15\] rf.registers\[29\]\[15\] rf.registers\[30\]\[15\]
+ rf.registers\[31\]\[15\] _1782_ _1680_ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4303_ _1025_ _1039_ _1058_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__o21ai_2
X_8071_ rf.registers\[20\]\[15\] _3487_ _4000_ VGND VGND VPWR VPWR _4006_ sky130_fd_sc_hd__mux2_1
X_5283_ _1171_ _1094_ _1098_ _1102_ _1109_ VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__a32oi_4
X_7022_ _3433_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4746__S _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8218__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5431__A _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8973_ clknet_leaf_40_clk _0133_ VGND VGND VPWR VPWR rf.registers\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6961__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7924_ net448 _3476_ _3927_ VGND VGND VPWR VPWR _3928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7855_ _3879_ VGND VGND VPWR VPWR _3891_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7358__A _3627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6806_ net993 _3120_ _3315_ VGND VGND VPWR VPWR _3319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_42_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7786_ _3854_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__clkbuf_1
X_4998_ _1671_ _1744_ _1749_ _1753_ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__o22a_1
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9525_ clknet_leaf_31_clk _0685_ VGND VGND VPWR VPWR rf.registers\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6737_ _3050_ net952 _3278_ VGND VGND VPWR VPWR _3282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7792__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6668_ _3245_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__clkbuf_1
X_9456_ clknet_leaf_7_clk _0616_ VGND VGND VPWR VPWR rf.registers\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_57_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5619_ _2255_ _2364_ _2371_ _2373_ VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__o211a_1
X_8407_ net139 _3483_ _4180_ VGND VGND VPWR VPWR _4184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9387_ clknet_leaf_4_clk _0547_ VGND VGND VPWR VPWR rf.registers\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6599_ _3048_ net553 _3206_ VGND VGND VPWR VPWR _3209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5606__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8338_ _4147_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5325__B _2080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8269_ _3118_ net227 _4108_ VGND VGND VPWR VPWR _4111_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5563__S0 _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4366__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6437__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7032__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7967__S _3915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5943__A1 _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5516__A _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4357__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4566__S _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7877__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6781__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5970_ _2140_ _2711_ VGND VGND VPWR VPWR _2712_ sky130_fd_sc_hd__xnor2_1
X_4921_ net2 VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__clkbuf_4
X_7640_ _3777_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
X_4852_ _1606_ _1607_ _1178_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7571_ _3031_ net1097 _3736_ VGND VGND VPWR VPWR _3741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4783_ rf.registers\[0\]\[9\] rf.registers\[1\]\[9\] rf.registers\[2\]\[9\] rf.registers\[3\]\[9\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4293__S0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9310_ clknet_leaf_73_clk _0470_ VGND VGND VPWR VPWR rf.registers\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6522_ net176 _3111_ _3157_ VGND VGND VPWR VPWR _3167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6453_ net20 VGND VGND VPWR VPWR _3124_ sky130_fd_sc_hd__buf_2
X_9241_ clknet_leaf_18_clk _0401_ VGND VGND VPWR VPWR rf.registers\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload40 clknet_leaf_63_clk VGND VGND VPWR VPWR clkload40/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__7117__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5404_ _1640_ _2151_ _2159_ VGND VGND VPWR VPWR _2160_ sky130_fd_sc_hd__o21a_2
Xclkload51 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload51/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4330__A _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload62 clknet_leaf_41_clk VGND VGND VPWR VPWR clkload62/Y sky130_fd_sc_hd__inv_8
X_9172_ clknet_leaf_29_clk _0332_ VGND VGND VPWR VPWR rf.registers\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6384_ _3076_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8123_ _4033_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5335_ rf.registers\[0\]\[1\] rf.registers\[1\]\[1\] rf.registers\[2\]\[1\] rf.registers\[3\]\[1\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2091_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5838__A1_N _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8054_ net537 _3470_ _3989_ VGND VGND VPWR VPWR _3997_ sky130_fd_sc_hd__mux2_1
X_5266_ rf.registers\[24\]\[24\] rf.registers\[25\]\[24\] rf.registers\[26\]\[24\]
+ rf.registers\[27\]\[24\] _1918_ _1919_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__mux4_1
XANTENNA__5545__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7005_ net178 _3113_ _3424_ VGND VGND VPWR VPWR _3425_ sky130_fd_sc_hd__mux2_1
X_5197_ _1901_ _1952_ _1766_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__a21o_1
XANTENNA__4673__A1 _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8956_ clknet_leaf_18_clk _0116_ VGND VGND VPWR VPWR rf.registers\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7907_ net217 _3460_ _3916_ VGND VGND VPWR VPWR _3919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8887_ clknet_leaf_33_clk _0047_ VGND VGND VPWR VPWR rf.registers\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7088__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7838_ _3882_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5100__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7769_ net333 _3458_ _3844_ VGND VGND VPWR VPWR _3846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_3_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_74_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9508_ clknet_leaf_62_clk _0668_ VGND VGND VPWR VPWR rf.registers\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8411__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9439_ clknet_leaf_73_clk _0599_ VGND VGND VPWR VPWR rf.registers\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4339__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4386__S _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6169__A1 _2613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4415__A _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5916__A1 _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4275__S0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold708 rf.registers\[5\]\[30\] VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold719 rf.registers\[28\]\[18\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5120_ _1860_ _1875_ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__nand2_1
XANTENNA__5527__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5051_ _1805_ _1806_ _1739_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8810_ clknet_leaf_6_clk _0994_ VGND VGND VPWR VPWR rf.registers\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8741_ clknet_leaf_61_clk _0925_ VGND VGND VPWR VPWR rf.registers\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5953_ _2340_ _2608_ _1879_ VGND VGND VPWR VPWR _2696_ sky130_fd_sc_hd__mux2_1
XANTENNA__4502__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4904_ _1640_ _1650_ _1654_ _1659_ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__a2bb2o_2
X_8672_ clknet_leaf_70_clk _0856_ VGND VGND VPWR VPWR rf.registers\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_5884_ net114 _1542_ VGND VGND VPWR VPWR _2630_ sky130_fd_sc_hd__or2b_1
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7623_ _3083_ net752 _3758_ VGND VGND VPWR VPWR _3768_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__9283__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4835_ rf.registers\[20\]\[17\] rf.registers\[21\]\[17\] rf.registers\[22\]\[17\]
+ rf.registers\[23\]\[17\] _1291_ _1194_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5907__B2 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4766_ rf.registers\[8\]\[8\] rf.registers\[9\]\[8\] rf.registers\[10\]\[8\] rf.registers\[11\]\[8\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__mux4_1
X_7554_ _3731_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6505_ _3158_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_60_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7485_ _3081_ net640 _3686_ VGND VGND VPWR VPWR _3695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4697_ rf.registers\[24\]\[12\] rf.registers\[25\]\[12\] rf.registers\[26\]\[12\]
+ rf.registers\[27\]\[12\] net100 _1221_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9224_ clknet_leaf_65_clk _0384_ VGND VGND VPWR VPWR rf.registers\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6436_ _3112_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6686__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9155_ clknet_leaf_53_clk _0315_ VGND VGND VPWR VPWR rf.registers\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6367_ _3022_ VGND VGND VPWR VPWR _3065_ sky130_fd_sc_hd__clkbuf_8
X_5318_ rf.registers\[12\]\[2\] rf.registers\[13\]\[2\] rf.registers\[14\]\[2\] rf.registers\[15\]\[2\]
+ _1673_ _1690_ VGND VGND VPWR VPWR _2074_ sky130_fd_sc_hd__mux4_1
X_8106_ _3155_ _3626_ VGND VGND VPWR VPWR _4024_ sky130_fd_sc_hd__nor2b_4
XANTENNA__5518__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9086_ clknet_leaf_74_clk _0246_ VGND VGND VPWR VPWR rf.registers\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6298_ net38 VGND VGND VPWR VPWR _3017_ sky130_fd_sc_hd__clkbuf_2
X_8037_ _3021_ VGND VGND VPWR VPWR _3987_ sky130_fd_sc_hd__inv_2
X_5249_ _2003_ _2004_ _1726_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__mux2_1
Xhold57 rf.registers\[12\]\[13\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 rf.registers\[1\]\[1\] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 rf.registers\[2\]\[12\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4741__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7596__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8939_ clknet_leaf_4_clk _0099_ VGND VGND VPWR VPWR rf.registers\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7348__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8141__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6450__A net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5066__A _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4980__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5005__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4732__S1 _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8316__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkload4_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4496__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ rf.registers\[4\]\[24\] rf.registers\[5\]\[24\] rf.registers\[6\]\[24\] rf.registers\[7\]\[24\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__mux4_1
XANTENNA__6360__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6562__A1 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4799__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4573__B1 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4551_ rf.registers\[12\]\[27\] rf.registers\[13\]\[27\] rf.registers\[14\]\[27\]
+ rf.registers\[15\]\[27\] net1164 _1268_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold505 rf.registers\[22\]\[8\] VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
X_7270_ _3071_ net812 _3577_ VGND VGND VPWR VPWR _3581_ sky130_fd_sc_hd__mux2_1
X_4482_ _1217_ _1237_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nand2_2
Xhold516 rf.registers\[10\]\[16\] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold527 rf.registers\[4\]\[10\] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 rf.registers\[3\]\[22\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _2421_ _2941_ _2943_ _2948_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__o22a_2
Xhold549 rf.registers\[16\]\[20\] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4420__S0 _1173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6152_ _2877_ _2879_ _2883_ VGND VGND VPWR VPWR _2884_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5103_ _1842_ _1858_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6083_ _2808_ _2818_ VGND VGND VPWR VPWR _2819_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_29_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5034_ rf.registers\[8\]\[20\] rf.registers\[9\]\[20\] rf.registers\[10\]\[20\] rf.registers\[11\]\[20\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_142_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8226__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7130__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6985_ _3414_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6250__B1 _1127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4487__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8724_ clknet_leaf_30_clk _0908_ VGND VGND VPWR VPWR rf.registers\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_5936_ _2486_ _2588_ _2679_ _1962_ _2333_ VGND VGND VPWR VPWR _2680_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_62_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8655_ clknet_leaf_28_clk _0839_ VGND VGND VPWR VPWR rf.registers\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5867_ _1087_ _2613_ VGND VGND VPWR VPWR _2614_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_38_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7606_ _3759_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4818_ rf.registers\[24\]\[16\] rf.registers\[25\]\[16\] rf.registers\[26\]\[16\]
+ rf.registers\[27\]\[16\] _1291_ _1194_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__mux4_1
X_8586_ clknet_leaf_8_clk _0770_ VGND VGND VPWR VPWR rf.registers\[22\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_5798_ _2499_ _2547_ _2347_ VGND VGND VPWR VPWR _2548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7537_ _3064_ net932 _3722_ VGND VGND VPWR VPWR _3723_ sky130_fd_sc_hd__mux2_1
X_4749_ _1503_ _1504_ _1190_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7468_ _3663_ VGND VGND VPWR VPWR _3686_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9207_ clknet_leaf_33_clk _0367_ VGND VGND VPWR VPWR rf.registers\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6419_ net40 VGND VGND VPWR VPWR _3101_ sky130_fd_sc_hd__buf_2
X_7399_ _3649_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5614__A _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8058__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput58 net58 VGND VGND VPWR VPWR alu_out[18] sky130_fd_sc_hd__buf_4
X_9138_ clknet_leaf_39_clk _0298_ VGND VGND VPWR VPWR rf.registers\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xoutput69 net69 VGND VGND VPWR VPWR alu_out[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_73_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9069_ clknet_leaf_40_clk _0229_ VGND VGND VPWR VPWR rf.registers\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4478__S0 _1182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7975__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7741__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4839__S _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4402__S0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4953__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4705__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5283__A1 _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8046__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4878__A1_N _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7885__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6232__B1 _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4469__S0 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5586__A2 _1874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6770_ _3083_ net1056 _3289_ VGND VGND VPWR VPWR _3299_ sky130_fd_sc_hd__mux2_1
XANTENNA__5130__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5721_ _2473_ _2385_ _1146_ VGND VGND VPWR VPWR _2474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6090__A _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8440_ net565 net35 _4191_ VGND VGND VPWR VPWR _4201_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5652_ _1666_ _2406_ VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__or2_1
XANTENNA__7732__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4603_ _1355_ _1358_ _1214_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__mux2_1
X_5583_ _1167_ _1661_ VGND VGND VPWR VPWR _2338_ sky130_fd_sc_hd__nor2_1
X_8371_ _4164_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4534_ _1065_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__buf_12
X_7322_ _3608_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_152_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4816__A1_N _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold302 rf.registers\[5\]\[17\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_152_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold313 rf.registers\[9\]\[14\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 rf.registers\[1\]\[11\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 rf.registers\[11\]\[0\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold346 rf.registers\[13\]\[9\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _1053_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__clkbuf_4
X_7253_ _3054_ net1145 _3566_ VGND VGND VPWR VPWR _3572_ sky130_fd_sc_hd__mux2_1
XANTENNA__4749__S _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold357 rf.registers\[24\]\[6\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold368 rf.registers\[8\]\[23\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 rf.registers\[21\]\[12\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
X_6204_ _1958_ _2931_ VGND VGND VPWR VPWR _2932_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7184_ _3534_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4396_ _1150_ _1151_ _1035_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6135_ _2847_ _2866_ _1147_ VGND VGND VPWR VPWR _2867_ sky130_fd_sc_hd__mux2_1
Xhold1002 rf.registers\[31\]\[26\] VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 rf.registers\[28\]\[15\] VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8460__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6066_ _2735_ _2801_ _2252_ VGND VGND VPWR VPWR _2802_ sky130_fd_sc_hd__mux2_1
Xhold1024 rf.registers\[25\]\[22\] VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 rf.registers\[14\]\[4\] VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 rf.registers\[20\]\[18\] VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ _1717_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__buf_4
Xhold1057 rf.registers\[21\]\[27\] VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 rf.registers\[23\]\[0\] VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__A_N _1528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6968_ _3404_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_46_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8707_ clknet_leaf_60_clk _0891_ VGND VGND VPWR VPWR rf.registers\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5919_ _2661_ _2662_ VGND VGND VPWR VPWR _2663_ sky130_fd_sc_hd__nand2_2
XFILLER_0_76_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6899_ net185 _3145_ _3362_ VGND VGND VPWR VPWR _3368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8638_ clknet_leaf_72_clk _0822_ VGND VGND VPWR VPWR rf.registers\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4537__B1 _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8569_ clknet_leaf_18_clk _0753_ VGND VGND VPWR VPWR rf.registers\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4632__S0 _1219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold880 rf.registers\[24\]\[25\] VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 rf.registers\[25\]\[2\] VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6874__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5998__B _2737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4871__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5254__A _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4926__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8442__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7940_ net191 _3493_ _3927_ VGND VGND VPWR VPWR _3936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5351__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7871_ _3899_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8504__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6822_ _3327_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4767__B1 _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9541_ clknet_leaf_61_clk _0701_ VGND VGND VPWR VPWR rf.registers\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6753_ _3290_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5704_ _2456_ VGND VGND VPWR VPWR _2457_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4333__A _1041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9472_ clknet_leaf_60_clk _0632_ VGND VGND VPWR VPWR rf.registers\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_154_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6684_ net758 _3134_ _3253_ VGND VGND VPWR VPWR _3254_ sky130_fd_sc_hd__mux2_1
X_8423_ _4192_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6959__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5635_ _2382_ _2389_ _2251_ VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__mux2_4
XFILLER_0_115_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7181__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4755__A1_N _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8354_ net631 _3497_ _4155_ VGND VGND VPWR VPWR _4156_ sky130_fd_sc_hd__mux2_1
X_5566_ _1696_ _2321_ _1670_ VGND VGND VPWR VPWR _2322_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold110 rf.registers\[11\]\[14\] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
X_7305_ _3599_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
Xhold121 rf.registers\[19\]\[6\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4479__S _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold132 rf.registers\[5\]\[12\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ rf.registers\[4\]\[21\] rf.registers\[5\]\[21\] rf.registers\[6\]\[21\] rf.registers\[7\]\[21\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5497_ _2179_ _2250_ _2252_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__mux2_1
X_8285_ _4096_ VGND VGND VPWR VPWR _4119_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_57_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold143 rf.registers\[4\]\[13\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold154 rf.registers\[19\]\[8\] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5615__A_N _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold165 rf.registers\[4\]\[3\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 rf.registers\[16\]\[0\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
X_7236_ _3037_ net512 _3555_ VGND VGND VPWR VPWR _3563_ sky130_fd_sc_hd__mux2_1
X_4448_ rf.registers\[8\]\[29\] rf.registers\[9\]\[29\] rf.registers\[10\]\[29\] rf.registers\[11\]\[29\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__mux4_1
Xhold187 rf.registers\[12\]\[5\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 rf.registers\[17\]\[18\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6694__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4379_ _1131_ _1134_ _1037_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__mux2_2
X_7167_ _3525_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _2408_ _2845_ _2846_ _2851_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__o22a_1
X_7098_ net18 VGND VGND VPWR VPWR _3483_ sky130_fd_sc_hd__buf_2
X_6049_ _1820_ _2768_ VGND VGND VPWR VPWR _2786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4942__S _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5030__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8424__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5238__A1 _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4418__A _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6986__A1 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5333__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4997__B1 _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4852__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8324__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6779__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5420_ _1758_ _2175_ _1800_ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5351_ rf.registers\[16\]\[15\] rf.registers\[17\]\[15\] rf.registers\[18\]\[15\]
+ rf.registers\[19\]\[15\] _1782_ _1680_ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4302_ _1046_ _1051_ _1056_ _1038_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8070_ _4005_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__clkbuf_1
X_5282_ _1962_ _2037_ _1879_ VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__mux2_4
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7021_ net438 _3130_ _3424_ VGND VGND VPWR VPWR _3433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7403__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4328__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8972_ clknet_leaf_49_clk _0132_ VGND VGND VPWR VPWR rf.registers\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_7923_ _3915_ VGND VGND VPWR VPWR _3927_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8234__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4762__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7854_ _3890_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5088__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6805_ _3318_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7785_ net233 _3474_ _3844_ VGND VGND VPWR VPWR _3854_ sky130_fd_sc_hd__mux2_1
X_4997_ _1717_ _1752_ _1729_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4835__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9524_ clknet_leaf_30_clk _0684_ VGND VGND VPWR VPWR rf.registers\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6736_ _3281_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9455_ clknet_leaf_28_clk _0615_ VGND VGND VPWR VPWR rf.registers\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6667_ net872 _3118_ _3242_ VGND VGND VPWR VPWR _3245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8406_ _4183_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5618_ _2372_ VGND VGND VPWR VPWR _2373_ sky130_fd_sc_hd__clkbuf_4
X_9386_ clknet_leaf_64_clk _0546_ VGND VGND VPWR VPWR rf.registers\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6598_ _3208_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8337_ net947 _3481_ _4144_ VGND VGND VPWR VPWR _4147_ sky130_fd_sc_hd__mux2_1
X_5549_ _1728_ _2296_ _2300_ _2304_ VGND VGND VPWR VPWR _2305_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_42_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8268_ _4110_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7219_ net13 net12 net11 VGND VGND VPWR VPWR _3553_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_6_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8409__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8199_ net406 _3479_ _4072_ VGND VGND VPWR VPWR _4074_ sky130_fd_sc_hd__mux2_1
XANTENNA__5563__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7313__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5622__A _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4672__S _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6453__A net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5079__S0 _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7983__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6599__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4701__A _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5251__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4903__B1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5008__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5003__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5532__A _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output52_A net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6959__A1 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8054__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4920_ _1675_ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__buf_4
XANTENNA__6363__A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4851_ rf.registers\[24\]\[19\] rf.registers\[25\]\[19\] rf.registers\[26\]\[19\]
+ rf.registers\[27\]\[19\] net127 _1222_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__mux4_1
XANTENNA__7893__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7570_ _3740_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4782_ rf.registers\[4\]\[9\] rf.registers\[5\]\[9\] rf.registers\[6\]\[9\] rf.registers\[7\]\[9\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__mux4_1
XANTENNA__4293__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6521_ _3166_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7136__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9240_ clknet_leaf_26_clk _0400_ VGND VGND VPWR VPWR rf.registers\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5147__B1 _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6452_ _3123_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload30 clknet_leaf_58_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__inv_8
XFILLER_0_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload41 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload41/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5403_ _2153_ _2155_ _2158_ net4 net5 VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__a221o_1
Xclkload52 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload52/Y sky130_fd_sc_hd__clkinv_4
X_9171_ clknet_leaf_32_clk _0331_ VGND VGND VPWR VPWR rf.registers\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4330__B _1085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload63 clknet_leaf_42_clk VGND VGND VPWR VPWR clkload63/Y sky130_fd_sc_hd__clkinvlp_4
X_6383_ _3075_ net1055 _3065_ VGND VGND VPWR VPWR _3076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8122_ net452 _3470_ _4025_ VGND VGND VPWR VPWR _4033_ sky130_fd_sc_hd__mux2_1
X_5334_ _1645_ _2089_ VGND VGND VPWR VPWR _2090_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8053_ _3996_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__clkbuf_1
X_5265_ rf.registers\[28\]\[24\] rf.registers\[29\]\[24\] rf.registers\[30\]\[24\]
+ rf.registers\[31\]\[24\] _1918_ _1919_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__mux4_1
XANTENNA__7133__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5545__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7004_ _3412_ VGND VGND VPWR VPWR _3424_ sky130_fd_sc_hd__clkbuf_8
X_5196_ rf.registers\[0\]\[28\] rf.registers\[1\]\[28\] rf.registers\[2\]\[28\] rf.registers\[3\]\[28\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__mux4_1
X_8955_ clknet_leaf_22_clk _0115_ VGND VGND VPWR VPWR rf.registers\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_7906_ _3918_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__clkbuf_1
X_8886_ clknet_leaf_24_clk _0046_ VGND VGND VPWR VPWR rf.registers\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7837_ _3095_ net1005 _3880_ VGND VGND VPWR VPWR _3882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4808__S0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7768_ _3845_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9507_ clknet_leaf_61_clk _0667_ VGND VGND VPWR VPWR rf.registers\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xclkload2 clknet_3_2__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
X_6719_ _3272_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7127__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7699_ _3019_ net1040 _3808_ VGND VGND VPWR VPWR _3809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7308__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5617__A _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9438_ clknet_leaf_71_clk _0598_ VGND VGND VPWR VPWR rf.registers\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5233__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9369_ clknet_leaf_22_clk _0529_ VGND VGND VPWR VPWR rf.registers\[20\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8139__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6882__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6183__A _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6169__A2 _2737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4275__S1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4431__A _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold709 rf.registers\[21\]\[8\] VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5527__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5050_ rf.registers\[16\]\[18\] rf.registers\[17\]\[18\] rf.registers\[18\]\[18\]
+ rf.registers\[19\]\[18\] _1719_ _1722_ VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8740_ clknet_leaf_62_clk _0924_ VGND VGND VPWR VPWR rf.registers\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5952_ _2503_ _2693_ _2694_ VGND VGND VPWR VPWR _2695_ sky130_fd_sc_hd__or3_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4903_ _1655_ _1658_ net5 VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__a21oi_1
X_8671_ clknet_leaf_73_clk _0855_ VGND VGND VPWR VPWR rf.registers\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5883_ _2427_ _2591_ _2628_ _2504_ VGND VGND VPWR VPWR _2629_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7622_ _3767_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4834_ rf.registers\[16\]\[17\] rf.registers\[17\]\[17\] rf.registers\[18\]\[17\]
+ rf.registers\[19\]\[17\] _1291_ _1194_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__mux4_1
XANTENNA__8512__S _4204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7553_ _3081_ net626 _3722_ VGND VGND VPWR VPWR _3731_ sky130_fd_sc_hd__mux2_1
X_4765_ _1107_ _1520_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6504_ net209 _3089_ _3157_ VGND VGND VPWR VPWR _3158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7484_ _3694_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4591__B2 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4696_ rf.registers\[28\]\[12\] rf.registers\[29\]\[12\] rf.registers\[30\]\[12\]
+ rf.registers\[31\]\[12\] net100 _1221_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__mux4_1
XANTENNA__5215__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9223_ clknet_leaf_66_clk _0383_ VGND VGND VPWR VPWR rf.registers\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6967__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6435_ net1003 _3111_ _3093_ VGND VGND VPWR VPWR _3112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9154_ clknet_leaf_55_clk _0314_ VGND VGND VPWR VPWR rf.registers\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6366_ net26 VGND VGND VPWR VPWR _3064_ sky130_fd_sc_hd__buf_2
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8105_ _4023_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__clkbuf_1
X_5317_ _1684_ _2072_ VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__and2_1
X_9085_ clknet_leaf_3_clk _0245_ VGND VGND VPWR VPWR rf.registers\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6268__A _1334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5518__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6297_ _3016_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__clkbuf_1
X_8036_ _3986_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__clkbuf_1
X_5248_ rf.registers\[24\]\[25\] rf.registers\[25\]\[25\] rf.registers\[26\]\[25\]
+ rf.registers\[27\]\[25\] _1822_ _1823_ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__mux4_1
XANTENNA__7798__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold58 rf.registers\[7\]\[11\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 rf.registers\[2\]\[4\] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _1889_ _1934_ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8938_ clknet_leaf_6_clk _0098_ VGND VGND VPWR VPWR rf.registers\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4516__A _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8869_ clknet_leaf_62_clk _0029_ VGND VGND VPWR VPWR rf.registers\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8422__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_rebuffer24_A _1298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7562__A _3735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7501__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5810__A _2286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4426__A net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4496__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5956__S _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4860__S _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6641__A _3230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6011__B2 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4573__A1 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4550_ _1302_ _1305_ _1187_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold506 rf.registers\[0\]\[25\] VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6787__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4481_ _1171_ _1228_ _1236_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a21oi_4
XANTENNA__5691__S _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold517 rf.registers\[10\]\[22\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold528 rf.registers\[9\]\[8\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ _1060_ _2678_ _2737_ _2947_ VGND VGND VPWR VPWR _2948_ sky130_fd_sc_hd__o22a_1
Xhold539 rf.registers\[19\]\[26\] VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4420__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6151_ _2812_ _2878_ _2882_ VGND VGND VPWR VPWR _2883_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6088__A _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5102_ _1672_ _1849_ _1853_ _1857_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__a2bb2o_2
X_6082_ _2812_ _2817_ VGND VGND VPWR VPWR _2818_ sky130_fd_sc_hd__nand2_1
XANTENNA__5825__A1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5825__B2 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5033_ _1785_ _1788_ _1699_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__mux2_1
XANTENNA__7411__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6984_ net715 _3089_ _3413_ VGND VGND VPWR VPWR _3414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6250__A1 _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4487__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8723_ clknet_leaf_34_clk _0907_ VGND VGND VPWR VPWR rf.registers\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5935_ _1666_ net81 _2251_ VGND VGND VPWR VPWR _2679_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4770__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8654_ clknet_leaf_44_clk _0838_ VGND VGND VPWR VPWR rf.registers\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_5866_ _2340_ _2487_ _2612_ _2530_ VGND VGND VPWR VPWR _2613_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_60_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7605_ _3064_ net1006 _3758_ VGND VGND VPWR VPWR _3759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4817_ _1528_ _1542_ _1558_ _1572_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__and4b_1
X_8585_ clknet_leaf_49_clk _0769_ VGND VGND VPWR VPWR rf.registers\[22\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5797_ _1669_ _2272_ _2325_ VGND VGND VPWR VPWR _2547_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7536_ _3699_ VGND VGND VPWR VPWR _3722_ sky130_fd_sc_hd__clkbuf_8
X_4748_ rf.registers\[12\]\[15\] rf.registers\[13\]\[15\] rf.registers\[14\]\[15\]
+ rf.registers\[15\]\[15\] _1201_ _1203_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7467_ _3685_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4679_ rf.registers\[24\]\[22\] rf.registers\[25\]\[22\] rf.registers\[26\]\[22\]
+ rf.registers\[27\]\[22\] _1182_ _1184_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9206_ clknet_leaf_24_clk _0366_ VGND VGND VPWR VPWR rf.registers\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6418_ _3100_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__clkbuf_1
X_7398_ _3062_ net856 _3639_ VGND VGND VPWR VPWR _3649_ sky130_fd_sc_hd__mux2_1
X_9137_ clknet_leaf_40_clk _0297_ VGND VGND VPWR VPWR rf.registers\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6349_ _3052_ net916 _3044_ VGND VGND VPWR VPWR _3053_ sky130_fd_sc_hd__mux2_1
Xoutput59 net59 VGND VGND VPWR VPWR alu_out[19] sky130_fd_sc_hd__buf_2
X_9068_ clknet_leaf_49_clk _0228_ VGND VGND VPWR VPWR rf.registers\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8019_ _3141_ net1154 _3974_ VGND VGND VPWR VPWR _3978_ sky130_fd_sc_hd__mux2_1
XANTENNA__8417__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7321__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clone44_A _1026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4478__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4680__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8152__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5427__S0 _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5201__C1 _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5077__A _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__9123__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4402__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5807__A1 _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4469__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5720_ _2381_ VGND VGND VPWR VPWR _2473_ sky130_fd_sc_hd__inv_2
XANTENNA__4590__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_44_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5651_ _2390_ _2405_ _2104_ VGND VGND VPWR VPWR _2406_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4602_ _1356_ _1357_ _1199_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8370_ net586 _3446_ _4155_ VGND VGND VPWR VPWR _4164_ sky130_fd_sc_hd__mux2_1
X_5582_ _2336_ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7321_ _3054_ net751 _3602_ VGND VGND VPWR VPWR _3608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4533_ _1287_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_152_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold303 rf.registers\[16\]\[31\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_152_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold314 rf.registers\[3\]\[28\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold325 rf.registers\[10\]\[26\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7252_ _3571_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
X_4464_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__buf_12
Xhold336 rf.registers\[6\]\[17\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 rf.registers\[12\]\[0\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold358 rf.registers\[17\]\[20\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 rf.registers\[9\]\[2\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ net98 _2930_ VGND VGND VPWR VPWR _2931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7183_ net394 _3487_ _3528_ VGND VGND VPWR VPWR _3534_ sky130_fd_sc_hd__mux2_1
X_4395_ rf.registers\[16\]\[0\] rf.registers\[17\]\[0\] rf.registers\[18\]\[0\] rf.registers\[19\]\[0\]
+ net94 _1061_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6134_ _1669_ _1732_ _2035_ VGND VGND VPWR VPWR _2866_ sky130_fd_sc_hd__a21oi_1
Xhold1003 rf.registers\[26\]\[9\] VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__dlygate4sd3_1
X_6065_ _2777_ _2800_ _1147_ VGND VGND VPWR VPWR _2801_ sky130_fd_sc_hd__mux2_1
Xhold1014 rf.registers\[0\]\[23\] VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 rf.registers\[15\]\[5\] VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 rf.registers\[21\]\[29\] VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 rf.registers\[19\]\[16\] VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8640__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5016_ _1766_ _1771_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__nand2_1
Xhold1058 rf.registers\[14\]\[21\] VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 rf.registers\[14\]\[16\] VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_37_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6967_ net616 _3145_ _3398_ VGND VGND VPWR VPWR _3404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8706_ clknet_leaf_60_clk _0890_ VGND VGND VPWR VPWR rf.registers\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5918_ _2175_ _2659_ _2660_ VGND VGND VPWR VPWR _2662_ sky130_fd_sc_hd__nand3_1
XFILLER_0_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4785__B2 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5982__B1 _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6898_ _3367_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_33_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__5409__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8637_ clknet_leaf_14_clk _0821_ VGND VGND VPWR VPWR rf.registers\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5849_ net115 _2596_ VGND VGND VPWR VPWR _2597_ sky130_fd_sc_hd__xor2_2
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4537__A1 _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8568_ clknet_leaf_21_clk _0752_ VGND VGND VPWR VPWR rf.registers\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4632__S1 _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7519_ _3713_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
X_8499_ _4232_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7487__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5625__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold870 rf.registers\[14\]\[13\] VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 rf.registers\[6\]\[30\] VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 rf.registers\[4\]\[7\] VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8147__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6456__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7051__S _3412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7411__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4871__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5725__B1 _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7226__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5489__C1 _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6366__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5270__A _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7870_ _3128_ net760 _3891_ VGND VGND VPWR VPWR _3899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6821_ net299 _3134_ _3326_ VGND VGND VPWR VPWR _3327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9540_ clknet_leaf_63_clk _0700_ VGND VGND VPWR VPWR rf.registers\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4767__A1 _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4311__S0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6752_ _3064_ net732 _3289_ VGND VGND VPWR VPWR _3290_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_15_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5703_ _2368_ _2367_ VGND VGND VPWR VPWR _2456_ sky130_fd_sc_hd__and2_1
X_9471_ clknet_leaf_71_clk _0631_ VGND VGND VPWR VPWR rf.registers\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_154_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6683_ _3230_ VGND VGND VPWR VPWR _3253_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_154_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8422_ net955 _3497_ _4191_ VGND VGND VPWR VPWR _4192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8520__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5634_ _2388_ VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5023__A1_N _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8353_ _4132_ VGND VGND VPWR VPWR _4155_ sky130_fd_sc_hd__clkbuf_8
X_5565_ _2319_ _2320_ _2044_ VGND VGND VPWR VPWR _2321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7136__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold100 rf.registers\[18\]\[1\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7469__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7304_ _3037_ net833 _3591_ VGND VGND VPWR VPWR _3599_ sky130_fd_sc_hd__mux2_1
Xhold111 rf.registers\[9\]\[30\] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _1214_ _1271_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__nand2_1
Xhold122 rf.registers\[6\]\[3\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
X_8284_ _4118_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__clkbuf_1
Xhold133 rf.registers\[17\]\[3\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ _2251_ VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold144 rf.registers\[5\]\[31\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
X_7235_ _3562_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
Xhold155 rf.registers\[19\]\[14\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6975__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4447_ _1202_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__buf_4
XFILLER_0_111_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold166 rf.registers\[18\]\[27\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold177 rf.registers\[19\]\[25\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 rf.registers\[3\]\[26\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 rf.registers\[19\]\[31\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7166_ net555 _3470_ _3517_ VGND VGND VPWR VPWR _3525_ sky130_fd_sc_hd__mux2_1
X_4378_ _1132_ _1133_ _1035_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _2549_ _2823_ _2731_ _2705_ _2850_ VGND VGND VPWR VPWR _2851_ sky130_fd_sc_hd__a221o_1
X_7097_ _3482_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
X_6048_ _1820_ _2768_ VGND VGND VPWR VPWR _2785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8197__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7999_ _3967_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8430__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6380__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5030__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6435__A1 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6914__A _3375_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4997__A1 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8188__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4434__A _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5964__S _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8360__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5350_ rf.registers\[20\]\[15\] rf.registers\[21\]\[15\] rf.registers\[22\]\[15\]
+ rf.registers\[23\]\[15\] _1734_ _1680_ VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4301_ net8 VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__buf_4
XANTENNA__6795__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5281_ _1999_ _2036_ _1877_ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__mux2_2
X_7020_ _3432_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_4_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__4685__B1 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4609__A _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4780__S0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6426__A1 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7623__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8971_ clknet_leaf_2_clk _0131_ VGND VGND VPWR VPWR rf.registers\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_7922_ _3926_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4532__S0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7853_ _3111_ net722 _3880_ VGND VGND VPWR VPWR _3890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7926__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6804_ net641 _3118_ _3315_ VGND VGND VPWR VPWR _3318_ sky130_fd_sc_hd__mux2_1
XANTENNA__5088__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7784_ _3853_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4996_ _1750_ _1751_ _1739_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__mux2_1
XANTENNA__4835__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6735_ _3048_ net312 _3278_ VGND VGND VPWR VPWR _3281_ sky130_fd_sc_hd__mux2_1
X_9523_ clknet_leaf_34_clk _0683_ VGND VGND VPWR VPWR rf.registers\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_83_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8250__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9454_ clknet_leaf_29_clk _0614_ VGND VGND VPWR VPWR rf.registers\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6666_ _3244_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8351__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5617_ _1060_ _2101_ VGND VGND VPWR VPWR _2372_ sky130_fd_sc_hd__and2_1
X_8405_ net885 _3481_ _4180_ VGND VGND VPWR VPWR _4183_ sky130_fd_sc_hd__mux2_1
X_9385_ clknet_leaf_50_clk _0545_ VGND VGND VPWR VPWR rf.registers\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6597_ _3046_ net239 _3206_ VGND VGND VPWR VPWR _3208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8336_ _4146_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5548_ _1696_ _2303_ _1670_ VGND VGND VPWR VPWR _2304_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8267_ _3116_ net527 _4108_ VGND VGND VPWR VPWR _4110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5479_ rf.registers\[16\]\[9\] rf.registers\[17\]\[9\] rf.registers\[18\]\[9\] rf.registers\[19\]\[9\]
+ _1675_ _1692_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__mux4_1
XANTENNA__6665__A1 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7862__A0 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5903__A _2567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7218_ net10 net9 net46 VGND VGND VPWR VPWR _3552_ sky130_fd_sc_hd__and3b_4
XTAP_TAPCELL_ROW_6_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8198_ _4073_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7149_ _3515_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5530__A1_N _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6417__A1 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7090__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7917__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5079__S1 _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8160__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5251__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4903__A1 _1655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7853__A0 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6656__A1 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5003__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7605__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4514__S0 net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8335__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4850_ rf.registers\[28\]\[19\] rf.registers\[29\]\[19\] rf.registers\[30\]\[19\]
+ rf.registers\[31\]\[19\] net127 _1222_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4781_ _1040_ _1536_ _1037_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__o21a_1
X_6520_ net297 _3109_ _3157_ VGND VGND VPWR VPWR _3166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8333__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6451_ net264 _3122_ _3114_ VGND VGND VPWR VPWR _3123_ sky130_fd_sc_hd__mux2_1
XANTENNA__5147__A1 _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload20 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__inv_8
XFILLER_0_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload31 clknet_leaf_59_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__clkinv_8
X_5402_ _2156_ _2157_ net3 VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload42 clknet_leaf_9_clk VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__clkinv_8
X_9170_ clknet_leaf_27_clk _0330_ VGND VGND VPWR VPWR rf.registers\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6382_ net31 VGND VGND VPWR VPWR _3075_ sky130_fd_sc_hd__clkbuf_2
Xclkload53 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload53/Y sky130_fd_sc_hd__inv_6
Xclkload64 clknet_leaf_43_clk VGND VGND VPWR VPWR clkload64/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8121_ _4032_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5333_ rf.registers\[4\]\[1\] rf.registers\[5\]\[1\] rf.registers\[6\]\[1\] rf.registers\[7\]\[1\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8052_ net723 _3468_ _3989_ VGND VGND VPWR VPWR _3996_ sky130_fd_sc_hd__mux2_1
X_5264_ _2018_ _2019_ _1901_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__mux2_1
XANTENNA__4658__B1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7003_ _3423_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5195_ _1889_ _1950_ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__and2_1
XANTENNA__4505__S0 _1220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8954_ clknet_leaf_17_clk _0114_ VGND VGND VPWR VPWR rf.registers\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7905_ net182 _3458_ _3916_ VGND VGND VPWR VPWR _3918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8885_ clknet_leaf_34_clk _0045_ VGND VGND VPWR VPWR rf.registers\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4830__B1 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7836_ _3881_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4808__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7767_ net183 _3454_ _3844_ VGND VGND VPWR VPWR _3845_ sky130_fd_sc_hd__mux2_1
X_4979_ _1721_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__buf_4
X_9506_ clknet_leaf_58_clk _0666_ VGND VGND VPWR VPWR rf.registers\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6718_ _3031_ net1117 _3267_ VGND VGND VPWR VPWR _3272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8324__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7698_ _3807_ VGND VGND VPWR VPWR _3808_ sky130_fd_sc_hd__clkbuf_8
Xclkload3 clknet_3_3__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinvlp_4
X_6649_ _3235_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__clkbuf_1
X_9437_ clknet_leaf_14_clk _0597_ VGND VGND VPWR VPWR rf.registers\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5233__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6886__A1 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9368_ clknet_leaf_27_clk _0528_ VGND VGND VPWR VPWR rf.registers\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8319_ _4137_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__clkbuf_1
X_9299_ clknet_leaf_37_clk _0459_ VGND VGND VPWR VPWR rf.registers\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4744__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7994__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7234__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4735__S0 net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8065__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5951_ _2522_ _2605_ _2591_ _2531_ VGND VGND VPWR VPWR _2694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4902_ _1656_ _1657_ _1645_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__mux2_1
X_8670_ clknet_leaf_72_clk _0854_ VGND VGND VPWR VPWR rf.registers\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5882_ _2441_ _2588_ _2590_ _2444_ VGND VGND VPWR VPWR _2628_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8554__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4833_ rf.registers\[28\]\[17\] rf.registers\[29\]\[17\] rf.registers\[30\]\[17\]
+ rf.registers\[31\]\[17\] _1191_ _1174_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__mux4_1
X_7621_ _3081_ net677 _3758_ VGND VGND VPWR VPWR _3767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7409__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7552_ _3730_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
X_4764_ rf.registers\[12\]\[8\] rf.registers\[13\]\[8\] rf.registers\[14\]\[8\] rf.registers\[15\]\[8\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6503_ _3156_ VGND VGND VPWR VPWR _3157_ sky130_fd_sc_hd__buf_4
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7483_ _3079_ net780 _3686_ VGND VGND VPWR VPWR _3694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4695_ _1449_ _1450_ _1036_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6868__A1 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5215__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9222_ clknet_leaf_66_clk _0382_ VGND VGND VPWR VPWR rf.registers\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6434_ net45 VGND VGND VPWR VPWR _3111_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9153_ clknet_leaf_57_clk _0313_ VGND VGND VPWR VPWR rf.registers\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6365_ _3063_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7144__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8104_ net251 _3452_ _3988_ VGND VGND VPWR VPWR _4023_ sky130_fd_sc_hd__mux2_1
X_5316_ rf.registers\[8\]\[2\] rf.registers\[9\]\[2\] rf.registers\[10\]\[2\] rf.registers\[11\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__mux4_1
X_9084_ clknet_leaf_16_clk _0244_ VGND VGND VPWR VPWR rf.registers\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6296_ net445 _3015_ _3007_ VGND VGND VPWR VPWR _3016_ sky130_fd_sc_hd__mux2_1
XANTENNA__6268__B _1904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8035_ _3017_ net826 _3951_ VGND VGND VPWR VPWR _3986_ sky130_fd_sc_hd__mux2_1
XANTENNA__4726__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5247_ rf.registers\[28\]\[25\] rf.registers\[29\]\[25\] rf.registers\[30\]\[25\]
+ rf.registers\[31\]\[25\] _1822_ _1823_ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__mux4_1
Xhold59 rf.registers\[9\]\[24\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ rf.registers\[4\]\[29\] rf.registers\[5\]\[29\] rf.registers\[6\]\[29\] rf.registers\[7\]\[29\]
+ _1767_ _1768_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__mux4_1
XANTENNA__7045__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8937_ clknet_leaf_47_clk _0097_ VGND VGND VPWR VPWR rf.registers\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5151__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8868_ clknet_leaf_48_clk _0028_ VGND VGND VPWR VPWR rf.registers\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7819_ net163 _3508_ _3866_ VGND VGND VPWR VPWR _3872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8799_ clknet_leaf_71_clk _0983_ VGND VGND VPWR VPWR rf.registers\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7319__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5628__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6859__A1 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_rebuffer17_A _1315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6459__A net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7054__S _3412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7989__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6893__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4717__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5390__S0 _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7036__A1 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6194__A _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4442__A _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4480_ _1230_ _1232_ _1205_ _1235_ _1215_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__o221a_4
Xhold507 rf.registers\[12\]\[28\] VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 rf.registers\[21\]\[17\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 rf.registers\[0\]\[19\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6150_ _2840_ _2843_ _2854_ _2880_ _2881_ VGND VGND VPWR VPWR _2882_ sky130_fd_sc_hd__o311a_1
XANTENNA__7899__S _3879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5101_ _1717_ _1856_ _1729_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__a21oi_1
X_6081_ _2814_ _2815_ _2748_ _2816_ VGND VGND VPWR VPWR _2817_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5032_ _1786_ _1787_ _1739_ VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__mux2_1
XANTENNA__5381__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5212__S _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6983_ _3412_ VGND VGND VPWR VPWR _3413_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8523__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8722_ clknet_leaf_27_clk _0906_ VGND VGND VPWR VPWR rf.registers\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5934_ _2502_ _2677_ _2104_ VGND VGND VPWR VPWR _2678_ sky130_fd_sc_hd__mux2_1
XANTENNA__8527__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5865_ _2426_ _2608_ _2611_ VGND VGND VPWR VPWR _2612_ sky130_fd_sc_hd__o21ai_1
X_8653_ clknet_leaf_43_clk _0837_ VGND VGND VPWR VPWR rf.registers\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4816_ _1025_ _1563_ _1567_ _1571_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__a2bb2o_4
X_7604_ _3735_ VGND VGND VPWR VPWR _3758_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8584_ clknet_leaf_49_clk _0768_ VGND VGND VPWR VPWR rf.registers\[22\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5796_ _2363_ _1758_ _2331_ _2419_ VGND VGND VPWR VPWR _2546_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4747_ rf.registers\[8\]\[15\] rf.registers\[9\]\[15\] rf.registers\[10\]\[15\] rf.registers\[11\]\[15\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__mux4_1
X_7535_ _3721_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
X_7466_ _3062_ net769 _3675_ VGND VGND VPWR VPWR _3685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4678_ rf.registers\[28\]\[22\] rf.registers\[29\]\[22\] rf.registers\[30\]\[22\]
+ rf.registers\[31\]\[22\] net135 _1184_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6417_ net215 _3099_ _3093_ VGND VGND VPWR VPWR _3100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9205_ clknet_leaf_31_clk _0365_ VGND VGND VPWR VPWR rf.registers\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_7397_ _3648_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput49 net49 VGND VGND VPWR VPWR alu_out[0] sky130_fd_sc_hd__buf_6
X_9136_ clknet_leaf_3_clk _0296_ VGND VGND VPWR VPWR rf.registers\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6348_ net19 VGND VGND VPWR VPWR _3052_ sky130_fd_sc_hd__clkbuf_2
X_9067_ clknet_leaf_4_clk _0227_ VGND VGND VPWR VPWR rf.registers\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6279_ net13 net11 net12 VGND VGND VPWR VPWR _3003_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_73_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7602__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8018_ _3977_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5372__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__9075__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8518__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5358__A _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5427__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_40_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_55_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4938__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5821__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5363__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4437__A _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5032__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6768__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5115__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8343__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5650_ _2404_ VGND VGND VPWR VPWR _2405_ sky130_fd_sc_hd__inv_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4601_ rf.registers\[24\]\[25\] rf.registers\[25\]\[25\] rf.registers\[26\]\[25\]
+ rf.registers\[27\]\[25\] _1351_ _1352_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__mux4_1
X_5581_ _1111_ _1126_ VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7320_ _3607_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4532_ rf.registers\[4\]\[26\] rf.registers\[5\]\[26\] rf.registers\[6\]\[26\] rf.registers\[7\]\[26\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_152_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold304 rf.registers\[7\]\[3\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 rf.registers\[28\]\[13\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
X_7251_ _3052_ net789 _3566_ VGND VGND VPWR VPWR _3571_ sky130_fd_sc_hd__mux2_1
Xhold326 rf.registers\[1\]\[2\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4463_ _1089_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__buf_12
XFILLER_0_13_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold337 rf.registers\[1\]\[20\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 rf.registers\[3\]\[29\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _2595_ _2929_ VGND VGND VPWR VPWR _2930_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold359 rf.registers\[30\]\[16\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7182_ _3533_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_4394_ rf.registers\[20\]\[0\] rf.registers\[21\]\[0\] rf.registers\[22\]\[0\] rf.registers\[23\]\[0\]
+ _1149_ _1061_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6133_ _2038_ _2864_ VGND VGND VPWR VPWR _2865_ sky130_fd_sc_hd__nor2_1
XANTENNA__8518__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1004 rf.registers\[15\]\[4\] VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__dlygate4sd3_1
X_6064_ _1840_ _1801_ VGND VGND VPWR VPWR _2800_ sky130_fd_sc_hd__and2b_1
Xhold1015 rf.registers\[28\]\[4\] VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5354__S0 _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1026 rf.registers\[26\]\[3\] VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__dlygate4sd3_1
X_5015_ _1769_ _1770_ _1713_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__mux2_1
Xhold1037 rf.registers\[26\]\[21\] VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 rf.registers\[27\]\[30\] VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1059 rf.registers\[29\]\[22\] VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5106__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6966_ _3403_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
X_8705_ clknet_leaf_61_clk _0889_ VGND VGND VPWR VPWR rf.registers\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5917_ _2660_ _2659_ _2175_ VGND VGND VPWR VPWR _2661_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6897_ net337 _3143_ _3362_ VGND VGND VPWR VPWR _3367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5409__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8636_ clknet_leaf_16_clk _0820_ VGND VGND VPWR VPWR rf.registers\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5848_ net121 _2593_ _2594_ _2595_ VGND VGND VPWR VPWR _2596_ sky130_fd_sc_hd__o31a_1
XFILLER_0_91_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8567_ _4267_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8489__A _4204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5779_ _1111_ VGND VGND VPWR VPWR _2530_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7518_ _3046_ net981 _3711_ VGND VGND VPWR VPWR _3713_ sky130_fd_sc_hd__mux2_1
X_8498_ net657 net30 _4227_ VGND VGND VPWR VPWR _4232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7449_ _3676_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold860 rf.registers\[18\]\[24\] VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 rf.registers\[16\]\[6\] VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 rf.registers\[29\]\[18\] VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 rf.registers\[27\]\[16\] VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9119_ clknet_leaf_74_clk _0279_ VGND VGND VPWR VPWR rf.registers\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8428__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7332__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6472__A net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7507__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6411__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output75_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5551__A _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_121_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6382__A net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8073__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6820_ _3303_ VGND VGND VPWR VPWR _3326_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4311__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6751_ _3266_ VGND VGND VPWR VPWR _3289_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5702_ _2339_ VGND VGND VPWR VPWR _2455_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9470_ clknet_leaf_73_clk _0630_ VGND VGND VPWR VPWR rf.registers\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6682_ _3252_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_154_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8421_ _4168_ VGND VGND VPWR VPWR _4191_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5633_ _2385_ _2387_ _1145_ VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7417__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5726__A _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6321__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5564_ rf.registers\[0\]\[5\] rf.registers\[1\]\[5\] rf.registers\[2\]\[5\] rf.registers\[3\]\[5\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2320_ sky130_fd_sc_hd__mux4_1
X_8352_ _4154_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_130_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold101 rf.registers\[9\]\[0\] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
X_7303_ _3598_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
X_4515_ _1269_ _1270_ _1190_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__mux2_1
Xhold112 rf.registers\[19\]\[3\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8283_ _3132_ net1131 _4108_ VGND VGND VPWR VPWR _4118_ sky130_fd_sc_hd__mux2_1
Xhold123 rf.registers\[19\]\[12\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ net86 VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__clkbuf_4
Xhold134 rf.registers\[24\]\[18\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold145 rf.registers\[13\]\[12\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
X_7234_ _3035_ net583 _3555_ VGND VGND VPWR VPWR _3562_ sky130_fd_sc_hd__mux2_1
X_4446_ _1029_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__clkbuf_4
Xhold156 rf.registers\[12\]\[31\] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 rf.registers\[12\]\[23\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 rf.registers\[7\]\[4\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold189 rf.registers\[29\]\[3\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8248__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7165_ _3524_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4377_ rf.registers\[24\]\[1\] rf.registers\[25\]\[1\] rf.registers\[26\]\[1\] rf.registers\[27\]\[1\]
+ net93 _1043_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__mux4_2
XANTENNA__7152__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6500__C_N net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _2495_ _2849_ _2503_ VGND VGND VPWR VPWR _2850_ sky130_fd_sc_hd__a21o_1
X_7096_ net321 _3481_ _3477_ VGND VGND VPWR VPWR _3482_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7641__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6047_ _1838_ _2783_ VGND VGND VPWR VPWR _2784_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6292__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7998_ _3120_ net614 _3963_ VGND VGND VPWR VPWR _3967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6949_ _3394_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8619_ clknet_leaf_5_clk _0803_ VGND VGND VPWR VPWR rf.registers\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7327__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5636__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8012__A _3951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8158__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5340__C1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold690 rf.registers\[14\]\[9\] VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7062__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5318__S0 _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5643__B1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7396__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6199__B2 _2737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4300_ _1054_ _1055_ _1047_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5280_ _2017_ _2035_ VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4685__A1 _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5309__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4780__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8970_ clknet_leaf_45_clk _0130_ VGND VGND VPWR VPWR rf.registers\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_7921_ net172 _3474_ _3916_ VGND VGND VPWR VPWR _3926_ sky130_fd_sc_hd__mux2_1
XANTENNA__4532__S1 _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7852_ _3889_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5220__S _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6803_ _3317_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7783_ net610 _3472_ _3844_ VGND VGND VPWR VPWR _3853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4995_ rf.registers\[0\]\[22\] rf.registers\[1\]\[22\] rf.registers\[2\]\[22\] rf.registers\[3\]\[22\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8531__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9522_ clknet_leaf_29_clk _0682_ VGND VGND VPWR VPWR rf.registers\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6734_ _3280_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9453_ clknet_leaf_8_clk _0613_ VGND VGND VPWR VPWR rf.registers\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6665_ net278 _3116_ _3242_ VGND VGND VPWR VPWR _3244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5456__A _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8404_ _4182_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5616_ _2366_ _2367_ _2370_ _2336_ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__a211o_1
X_9384_ clknet_leaf_49_clk _0544_ VGND VGND VPWR VPWR rf.registers\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6596_ _3207_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6986__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8335_ net788 _3479_ _4144_ VGND VGND VPWR VPWR _4146_ sky130_fd_sc_hd__mux2_1
X_5547_ _2301_ _2302_ _1738_ VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__mux2_1
XANTENNA__7311__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5478_ rf.registers\[20\]\[9\] rf.registers\[21\]\[9\] rf.registers\[22\]\[9\] rf.registers\[23\]\[9\]
+ _1675_ _1692_ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__mux4_1
X_8266_ _4109_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__clkbuf_1
X_7217_ _3551_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
X_4429_ rf.registers\[24\]\[29\] rf.registers\[25\]\[29\] rf.registers\[26\]\[29\]
+ rf.registers\[27\]\[29\] _1182_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__mux4_2
X_8197_ net920 _3476_ _4072_ VGND VGND VPWR VPWR _4073_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7148_ net866 _3452_ _3455_ VGND VGND VPWR VPWR _3515_ sky130_fd_sc_hd__mux2_1
X_7079_ net43 VGND VGND VPWR VPWR _3470_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4535__A _1290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4364__B1 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7520__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4514__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4445__A _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5040__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8351__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4780_ rf.registers\[12\]\[9\] rf.registers\[13\]\[9\] rf.registers\[14\]\[9\] rf.registers\[15\]\[9\]
+ net107 _1105_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6450_ net19 VGND VGND VPWR VPWR _3122_ sky130_fd_sc_hd__buf_2
Xclkload10 clknet_leaf_69_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__inv_8
Xclkload21 clknet_leaf_7_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_113_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload32 clknet_leaf_61_clk VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__clkinv_4
X_5401_ rf.registers\[12\]\[13\] rf.registers\[13\]\[13\] rf.registers\[14\]\[13\]
+ rf.registers\[15\]\[13\] _1702_ _1678_ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6381_ _3074_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__clkbuf_1
Xclkload43 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload43/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload54 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload54/Y sky130_fd_sc_hd__inv_6
Xclkload65 clknet_leaf_44_clk VGND VGND VPWR VPWR clkload65/Y sky130_fd_sc_hd__inv_6
XFILLER_0_101_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5332_ _2084_ _2085_ _2086_ _2087_ net3 _1655_ VGND VGND VPWR VPWR _2088_ sky130_fd_sc_hd__mux4_2
X_8120_ net439 _3468_ _4025_ VGND VGND VPWR VPWR _4032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8051_ _3995_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__clkbuf_1
X_5263_ rf.registers\[16\]\[24\] rf.registers\[17\]\[24\] rf.registers\[18\]\[24\]
+ rf.registers\[19\]\[24\] _1918_ _1919_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_149_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4658__A1 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7002_ net559 _3111_ _3413_ VGND VGND VPWR VPWR _3423_ sky130_fd_sc_hd__mux2_1
X_5194_ rf.registers\[4\]\[28\] rf.registers\[5\]\[28\] rf.registers\[6\]\[28\] rf.registers\[7\]\[28\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__mux4_1
X_8953_ clknet_leaf_19_clk _0113_ VGND VGND VPWR VPWR rf.registers\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4505__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7904_ _3917_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4355__A _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8884_ clknet_leaf_38_clk _0044_ VGND VGND VPWR VPWR rf.registers\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4830__A1 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7835_ _3089_ net1150 _3880_ VGND VGND VPWR VPWR _3881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7766_ _3843_ VGND VGND VPWR VPWR _3844_ sky130_fd_sc_hd__buf_4
X_4978_ _1733_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__clkbuf_8
X_9505_ clknet_leaf_57_clk _0665_ VGND VGND VPWR VPWR rf.registers\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6717_ _3271_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7697_ _3020_ _3553_ VGND VGND VPWR VPWR _3807_ sky130_fd_sc_hd__nand2_4
XFILLER_0_117_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload4 clknet_3_5__leaf_clk VGND VGND VPWR VPWR clkload4/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9436_ clknet_leaf_18_clk _0596_ VGND VGND VPWR VPWR rf.registers\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6648_ net579 _3099_ _3231_ VGND VGND VPWR VPWR _3235_ sky130_fd_sc_hd__mux2_1
XANTENNA__7532__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9367_ clknet_leaf_33_clk _0527_ VGND VGND VPWR VPWR rf.registers\[20\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6579_ _3198_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7605__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8088__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8318_ net398 _3462_ _4133_ VGND VGND VPWR VPWR _4137_ sky130_fd_sc_hd__mux2_1
X_9298_ clknet_leaf_37_clk _0458_ VGND VGND VPWR VPWR rf.registers\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8249_ _4100_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4744__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8436__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7340__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5782__C1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8079__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4735__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5950_ _2692_ _2679_ VGND VGND VPWR VPWR _2693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4901_ rf.registers\[0\]\[0\] rf.registers\[1\]\[0\] rf.registers\[2\]\[0\] rf.registers\[3\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5881_ _2335_ _2626_ VGND VGND VPWR VPWR _2627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7620_ _3766_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__clkbuf_1
X_4832_ rf.registers\[24\]\[17\] rf.registers\[25\]\[17\] rf.registers\[26\]\[17\]
+ rf.registers\[27\]\[17\] _1291_ _1194_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_47_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7551_ _3079_ net1062 _3722_ VGND VGND VPWR VPWR _3730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4763_ _1515_ _1518_ _1037_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__mux2_4
XFILLER_0_83_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4671__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6502_ _3153_ _3155_ VGND VGND VPWR VPWR _3156_ sky130_fd_sc_hd__nor2_4
X_4694_ rf.registers\[16\]\[12\] rf.registers\[17\]\[12\] rf.registers\[18\]\[12\]
+ rf.registers\[19\]\[12\] net100 _1221_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__mux4_1
X_7482_ _3693_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_60_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9221_ clknet_leaf_61_clk _0381_ VGND VGND VPWR VPWR rf.registers\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6433_ _3110_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9152_ clknet_leaf_68_clk _0312_ VGND VGND VPWR VPWR rf.registers\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6364_ _3062_ net719 _3044_ VGND VGND VPWR VPWR _3063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8103_ _4022_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__clkbuf_1
X_5315_ _2067_ _2070_ net4 VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__mux2_1
X_6295_ net37 VGND VGND VPWR VPWR _3015_ sky130_fd_sc_hd__clkbuf_2
X_9083_ clknet_leaf_36_clk _0243_ VGND VGND VPWR VPWR rf.registers\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_8034_ _3985_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8490__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5246_ _2000_ _2001_ _1726_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__mux2_1
XANTENNA__4726__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4784__S _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4500__B1 _1255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8256__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5177_ _1929_ _1932_ _1700_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__mux2_1
XANTENNA__7160__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8936_ clknet_leaf_63_clk _0096_ VGND VGND VPWR VPWR rf.registers\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5151__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8867_ clknet_leaf_68_clk _0027_ VGND VGND VPWR VPWR rf.registers\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6504__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7818_ _3871_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6556__A1 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8798_ clknet_leaf_0_clk _0982_ VGND VGND VPWR VPWR rf.registers\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7749_ _3073_ net980 _3830_ VGND VGND VPWR VPWR _3835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4662__S0 _1267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9419_ clknet_leaf_7_clk _0579_ VGND VGND VPWR VPWR rf.registers\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5819__A0 _2458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8481__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4717__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6475__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8166__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5390__S1 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7992__A0 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6414__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4558__B1 _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4869__S _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7245__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold508 rf.registers\[6\]\[22\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold519 rf.registers\[22\]\[31\] VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5100_ _1854_ _1855_ _1726_ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6080_ _2770_ _2809_ VGND VGND VPWR VPWR _2816_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5031_ rf.registers\[24\]\[20\] rf.registers\[25\]\[20\] rf.registers\[26\]\[20\]
+ rf.registers\[27\]\[20\] _1782_ _1680_ VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__mux4_1
XANTENNA__6385__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5381__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8224__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7983__A0 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6982_ _3090_ _3411_ VGND VGND VPWR VPWR _3412_ sky130_fd_sc_hd__nor2_4
XFILLER_0_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8721_ clknet_leaf_30_clk _0905_ VGND VGND VPWR VPWR rf.registers\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5933_ _2673_ _2676_ _2501_ VGND VGND VPWR VPWR _2677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4892__S0 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6324__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8652_ clknet_leaf_46_clk _0836_ VGND VGND VPWR VPWR rf.registers\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5864_ _2252_ _2610_ VGND VGND VPWR VPWR _2611_ sky130_fd_sc_hd__nand2_1
X_7603_ _3757_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_32_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4815_ _1088_ _1570_ net8 VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__a21oi_2
X_8583_ clknet_leaf_66_clk _0767_ VGND VGND VPWR VPWR rf.registers\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5795_ _2539_ _2540_ _2543_ VGND VGND VPWR VPWR _2545_ sky130_fd_sc_hd__or3_1
XANTENNA__4644__S0 _1104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7944__A _3915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7534_ _3062_ net976 _3711_ VGND VGND VPWR VPWR _3721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4746_ _1498_ _1501_ _1187_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7465_ _3684_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_1
X_4677_ _1431_ _1432_ _1178_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__mux2_1
X_9204_ clknet_leaf_42_clk _0364_ VGND VGND VPWR VPWR rf.registers\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6416_ net39 VGND VGND VPWR VPWR _3099_ sky130_fd_sc_hd__buf_2
X_7396_ _3060_ net266 _3639_ VGND VGND VPWR VPWR _3648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6994__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9135_ clknet_leaf_8_clk _0295_ VGND VGND VPWR VPWR rf.registers\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6347_ _3051_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__clkbuf_1
X_9066_ clknet_leaf_8_clk _0226_ VGND VGND VPWR VPWR rf.registers\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6278_ net32 VGND VGND VPWR VPWR _3002_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__5277__A1 _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8017_ _3139_ net734 _3974_ VGND VGND VPWR VPWR _3977_ sky130_fd_sc_hd__mux2_1
XANTENNA__6295__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5229_ rf.registers\[24\]\[26\] rf.registers\[25\]\[26\] rf.registers\[26\]\[26\]
+ rf.registers\[27\]\[26\] _1881_ _1883_ VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__mux4_1
XANTENNA__5372__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8215__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8919_ clknet_leaf_23_clk _0079_ VGND VGND VPWR VPWR rf.registers\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5639__A _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4543__A _1298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4635__S0 _1290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5201__B2 _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7065__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4938__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5060__S0 _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8454__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5821__B _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5363__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5115__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap81 _2039_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4874__S0 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4600_ rf.registers\[28\]\[25\] rf.registers\[29\]\[25\] rf.registers\[30\]\[25\]
+ rf.registers\[31\]\[25\] _1351_ _1352_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5580_ _1060_ _1085_ VGND VGND VPWR VPWR _2335_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4599__S _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4531_ _1048_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5284__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold305 rf.registers\[13\]\[3\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 rf.registers\[16\]\[3\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7250_ _3570_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4462_ rf.registers\[20\]\[28\] rf.registers\[21\]\[28\] rf.registers\[22\]\[28\]
+ rf.registers\[23\]\[28\] _1182_ _1184_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__mux4_2
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold327 rf.registers\[7\]\[14\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold338 rf.registers\[17\]\[21\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold349 rf.registers\[22\]\[13\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _1316_ _1385_ _2872_ VGND VGND VPWR VPWR _2929_ sky130_fd_sc_hd__or3_1
XANTENNA__4703__B1 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4393_ A2[0] VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__buf_12
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7181_ net409 _3485_ _3528_ VGND VGND VPWR VPWR _3533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7703__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6132_ _2104_ _2373_ VGND VGND VPWR VPWR _2864_ sky130_fd_sc_hd__nand2_1
X_6063_ _2583_ _2733_ _2426_ VGND VGND VPWR VPWR _2799_ sky130_fd_sc_hd__mux2_1
Xhold1005 rf.registers\[13\]\[26\] VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5354__S1 _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1016 rf.registers\[28\]\[27\] VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7004__A _3412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1027 rf.registers\[13\]\[15\] VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 rf.registers\[22\]\[22\] VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__dlygate4sd3_1
X_5014_ rf.registers\[12\]\[21\] rf.registers\[13\]\[21\] rf.registers\[14\]\[21\]
+ rf.registers\[15\]\[21\] _1767_ _1768_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__mux4_1
Xhold1049 rf.registers\[13\]\[19\] VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_37_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5106__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6965_ net937 _3143_ _3398_ VGND VGND VPWR VPWR _3403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8704_ clknet_leaf_69_clk _0888_ VGND VGND VPWR VPWR rf.registers\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_5916_ _2536_ _2658_ net1159 VGND VGND VPWR VPWR _2660_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6896_ _3366_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8635_ clknet_leaf_34_clk _0819_ VGND VGND VPWR VPWR rf.registers\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_5847_ net47 _2503_ VGND VGND VPWR VPWR _2595_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8566_ net887 net31 _3006_ VGND VGND VPWR VPWR _4267_ sky130_fd_sc_hd__mux2_1
X_5778_ _1666_ _2523_ _2528_ _2495_ VGND VGND VPWR VPWR _2529_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_134_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5290__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7517_ _3712_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__clkbuf_1
X_4729_ _1481_ _1482_ _1483_ _1484_ _1189_ _1078_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8497_ _4231_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7448_ _3043_ net889 _3675_ VGND VGND VPWR VPWR _3676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold850 rf.registers\[27\]\[20\] VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 rf.registers\[3\]\[11\] VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__dlygate4sd3_1
X_7379_ _3627_ VGND VGND VPWR VPWR _3639_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__7613__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold872 rf.registers\[25\]\[9\] VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__dlygate4sd3_1
X_9118_ clknet_leaf_74_clk _0278_ VGND VGND VPWR VPWR rf.registers\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold883 rf.registers\[20\]\[29\] VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 rf.registers\[27\]\[19\] VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__dlygate4sd3_1
X_9049_ clknet_leaf_19_clk _0209_ VGND VGND VPWR VPWR rf.registers\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6998__A1 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8444__S _4168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4856__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4273__A _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6899__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7175__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5186__B1 _1941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5725__A2 _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5489__A1 _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output68_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5978__S _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8354__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5279__A _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4847__S0 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6750_ _3288_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5701_ _2422_ _2436_ _2446_ _2454_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__o31a_4
XANTENNA__7166__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6681_ net939 _3132_ _3242_ VGND VGND VPWR VPWR _3252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7494__A _3699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8420_ _4190_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5632_ _1168_ _1997_ _2386_ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_116_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8351_ net421 _3495_ _4144_ VGND VGND VPWR VPWR _4154_ sky130_fd_sc_hd__mux2_1
X_5563_ rf.registers\[4\]\[5\] rf.registers\[5\]\[5\] rf.registers\[6\]\[5\] rf.registers\[7\]\[5\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2319_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7302_ _3035_ net750 _3591_ VGND VGND VPWR VPWR _3598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4514_ rf.registers\[12\]\[21\] rf.registers\[13\]\[21\] rf.registers\[14\]\[21\]
+ rf.registers\[15\]\[21\] net1164 _1268_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__mux4_1
X_8282_ _4117_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__clkbuf_1
Xhold102 rf.registers\[3\]\[20\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5494_ _2213_ _2249_ _2178_ VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__mux2_1
Xhold113 rf.registers\[1\]\[28\] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 rf.registers\[9\]\[17\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 rf.registers\[18\]\[2\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
X_7233_ _3561_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8529__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold146 rf.registers\[2\]\[11\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _1200_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__buf_12
Xhold157 rf.registers\[15\]\[11\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 rf.registers\[17\]\[4\] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7433__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold179 rf.registers\[1\]\[0\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7164_ net167 _3468_ _3517_ VGND VGND VPWR VPWR _3524_ sky130_fd_sc_hd__mux2_1
X_4376_ rf.registers\[28\]\[1\] rf.registers\[29\]\[1\] rf.registers\[30\]\[1\] rf.registers\[31\]\[1\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux4_2
X_6115_ _2778_ _2848_ _1879_ VGND VGND VPWR VPWR _2849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ net17 VGND VGND VPWR VPWR _3481_ sky130_fd_sc_hd__buf_2
XANTENNA__5101__B1 _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6046_ _1618_ _2782_ VGND VGND VPWR VPWR _2783_ sky130_fd_sc_hd__xor2_1
XANTENNA__4792__S _1034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6573__A _3194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5404__A1 _1640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7997_ _3966_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4838__S0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6948_ net468 _3126_ _3387_ VGND VGND VPWR VPWR _3394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6879_ _3357_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6512__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8618_ clknet_leaf_64_clk _0802_ VGND VGND VPWR VPWR rf.registers\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5263__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8549_ _4258_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_20_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8409__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold680 rf.registers\[31\]\[0\] VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold691 rf.registers\[21\]\[21\] VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4268__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5318__S1 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5643__A1 _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6199__A2 _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7518__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4731__A _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5006__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8349__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7253__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5562__A _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5309__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7920_ _3925_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8084__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4906__A _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7851_ _3109_ net929 _3880_ VGND VGND VPWR VPWR _3889_ sky130_fd_sc_hd__mux2_1
X_6802_ net501 _3116_ _3315_ VGND VGND VPWR VPWR _3317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7782_ _3852_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5937__A2 _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4994_ rf.registers\[4\]\[22\] rf.registers\[5\]\[22\] rf.registers\[6\]\[22\] rf.registers\[7\]\[22\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__mux4_1
X_9521_ clknet_leaf_29_clk _0681_ VGND VGND VPWR VPWR rf.registers\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6733_ _3046_ net174 _3278_ VGND VGND VPWR VPWR _3280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9452_ clknet_leaf_45_clk _0612_ VGND VGND VPWR VPWR rf.registers\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6664_ _3243_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5245__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8403_ net743 _3479_ _4180_ VGND VGND VPWR VPWR _4182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5615_ _2363_ _2368_ _2369_ VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__and3b_1
X_9383_ clknet_leaf_65_clk _0543_ VGND VGND VPWR VPWR rf.registers\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6595_ _3043_ net935 _3206_ VGND VGND VPWR VPWR _3207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8334_ _4145_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5546_ rf.registers\[0\]\[4\] rf.registers\[1\]\[4\] rf.registers\[2\]\[4\] rf.registers\[3\]\[4\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8265_ _3113_ net368 _4108_ VGND VGND VPWR VPWR _4109_ sky130_fd_sc_hd__mux2_1
X_5477_ _2231_ _2232_ _1712_ VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__mux2_1
X_7216_ net304 _3452_ _3516_ VGND VGND VPWR VPWR _3551_ sky130_fd_sc_hd__mux2_1
X_4428_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__buf_4
X_8196_ _4060_ VGND VGND VPWR VPWR _4072_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7147_ _3514_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_4359_ rf.registers\[20\]\[2\] rf.registers\[21\]\[2\] rf.registers\[22\]\[2\] rf.registers\[23\]\[2\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__mux4_2
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7078_ _3469_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
X_6029_ _1512_ _1602_ _2658_ _2536_ VGND VGND VPWR VPWR _2767_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_87_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5997__B_N _1085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7338__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6242__S _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4364__A1 _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6478__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_8_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6417__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5475__S0 _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload11 clknet_leaf_70_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__clkinv_8
X_5400_ rf.registers\[8\]\[13\] rf.registers\[9\]\[13\] rf.registers\[10\]\[13\] rf.registers\[11\]\[13\]
+ _1702_ _1678_ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload22 clknet_leaf_64_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__clkinv_4
Xclkload33 clknet_leaf_45_clk VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_113_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6380_ _3073_ net1064 _3065_ VGND VGND VPWR VPWR _3074_ sky130_fd_sc_hd__mux2_1
Xclkload44 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload44/Y sky130_fd_sc_hd__clkinv_8
Xclkload55 clknet_leaf_21_clk VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__inv_12
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5331_ rf.registers\[20\]\[1\] rf.registers\[21\]\[1\] rf.registers\[22\]\[1\] rf.registers\[23\]\[1\]
+ _1673_ _1690_ VGND VGND VPWR VPWR _2087_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload66 clknet_leaf_30_clk VGND VGND VPWR VPWR clkload66/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__8079__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8050_ net526 _3466_ _3989_ VGND VGND VPWR VPWR _3995_ sky130_fd_sc_hd__mux2_1
XANTENNA__4400__S _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5262_ rf.registers\[20\]\[24\] rf.registers\[21\]\[24\] rf.registers\[22\]\[24\]
+ rf.registers\[23\]\[24\] _1918_ _1919_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_149_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7001_ _3422_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
X_5193_ _1945_ _1946_ _1947_ _1948_ _1889_ _1773_ VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__mux4_1
XANTENNA__7711__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6327__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4636__A _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8952_ clknet_leaf_26_clk _0112_ VGND VGND VPWR VPWR rf.registers\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5231__S _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7903_ net662 _3454_ _3916_ VGND VGND VPWR VPWR _3917_ sky130_fd_sc_hd__mux2_1
X_8883_ clknet_leaf_36_clk _0043_ VGND VGND VPWR VPWR rf.registers\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_7834_ _3879_ VGND VGND VPWR VPWR _3880_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5466__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7765_ _3003_ _3091_ VGND VGND VPWR VPWR _3843_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_82_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4977_ _1702_ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__buf_4
XANTENNA__7158__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6716_ _3029_ net1031 _3267_ VGND VGND VPWR VPWR _3271_ sky130_fd_sc_hd__mux2_1
X_9504_ clknet_leaf_69_clk _0664_ VGND VGND VPWR VPWR rf.registers\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4371__A _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7696_ _3806_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5218__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload5 clknet_3_6__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_8
X_9435_ clknet_leaf_23_clk _0595_ VGND VGND VPWR VPWR rf.registers\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6647_ _3234_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9366_ clknet_leaf_24_clk _0526_ VGND VGND VPWR VPWR rf.registers\[20\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6578_ _3027_ net495 _3195_ VGND VGND VPWR VPWR _3198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8317_ _4136_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__clkbuf_1
X_5529_ _1828_ _2284_ _1728_ VGND VGND VPWR VPWR _2285_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9297_ clknet_leaf_41_clk _0457_ VGND VGND VPWR VPWR rf.registers\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6298__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8248_ _3097_ net848 _4097_ VGND VGND VPWR VPWR _4100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8179_ _4063_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7621__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8452__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7068__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6700__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6001__A _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5840__A _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output50_A net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5051__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4900_ rf.registers\[4\]\[0\] rf.registers\[5\]\[0\] rf.registers\[6\]\[0\] rf.registers\[7\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__mux4_1
XANTENNA__4890__S _1645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8362__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5880_ _2546_ _2570_ _2625_ _2105_ VGND VGND VPWR VPWR _2626_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_72_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4831_ _1215_ _1578_ _1582_ _1586_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7550_ _3729_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4762_ _1516_ _1517_ _1035_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6501_ _3154_ VGND VGND VPWR VPWR _3155_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4671__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7481_ _3077_ net229 _3686_ VGND VGND VPWR VPWR _3693_ sky130_fd_sc_hd__mux2_1
X_4693_ rf.registers\[20\]\[12\] rf.registers\[21\]\[12\] rf.registers\[22\]\[12\]
+ rf.registers\[23\]\[12\] net100 _1221_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9220_ clknet_leaf_63_clk _0380_ VGND VGND VPWR VPWR rf.registers\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6432_ net320 _3109_ _3093_ VGND VGND VPWR VPWR _3110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9151_ clknet_leaf_71_clk _0311_ VGND VGND VPWR VPWR rf.registers\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6363_ net24 VGND VGND VPWR VPWR _3062_ sky130_fd_sc_hd__clkbuf_2
X_8102_ net1099 _3450_ _3988_ VGND VGND VPWR VPWR _4022_ sky130_fd_sc_hd__mux2_1
X_5314_ _2068_ _2069_ _1645_ VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__mux2_1
X_9082_ clknet_leaf_37_clk _0242_ VGND VGND VPWR VPWR rf.registers\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6294_ _3014_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5828__A1 _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8033_ _3015_ net546 _3951_ VGND VGND VPWR VPWR _3985_ sky130_fd_sc_hd__mux2_1
XANTENNA__8537__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5245_ rf.registers\[16\]\[25\] rf.registers\[17\]\[25\] rf.registers\[18\]\[25\]
+ rf.registers\[19\]\[25\] _1822_ _1823_ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__mux4_1
XANTENNA__6846__A _3339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7441__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5176_ _1930_ _1931_ _1726_ VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__mux2_1
XANTENNA__7450__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6253__A1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8935_ clknet_leaf_2_clk _0095_ VGND VGND VPWR VPWR rf.registers\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8866_ clknet_leaf_56_clk _0026_ VGND VGND VPWR VPWR rf.registers\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_63_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5439__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7817_ net141 _3506_ _3866_ VGND VGND VPWR VPWR _3871_ sky130_fd_sc_hd__mux2_1
X_8797_ clknet_leaf_15_clk _0981_ VGND VGND VPWR VPWR rf.registers\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7748_ _3834_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4662__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7679_ net554 _3504_ _3794_ VGND VGND VPWR VPWR _3798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6520__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9418_ clknet_leaf_8_clk _0578_ VGND VGND VPWR VPWR rf.registers\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9349_ clknet_leaf_52_clk _0509_ VGND VGND VPWR VPWR rf.registers\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_95_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5819__A1 _2567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8182__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4350__S0 _1104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4558__A1 _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7526__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold509 rf.registers\[19\]\[7\] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7261__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5030_ rf.registers\[28\]\[20\] rf.registers\[29\]\[20\] rf.registers\[30\]\[20\]
+ rf.registers\[31\]\[20\] _1782_ _1680_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__mux4_1
XANTENNA__4494__B1 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ net10 net9 net46 VGND VGND VPWR VPWR _3411_ sky130_fd_sc_hd__nand3_4
XANTENNA__8092__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5932_ _2674_ _2675_ _1147_ VGND VGND VPWR VPWR _2676_ sky130_fd_sc_hd__mux2_1
XANTENNA__6605__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8720_ clknet_leaf_9_clk _0904_ VGND VGND VPWR VPWR rf.registers\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4914__A _1640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8651_ clknet_leaf_7_clk _0835_ VGND VGND VPWR VPWR rf.registers\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5863_ _2565_ _2609_ _1803_ VGND VGND VPWR VPWR _2610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7602_ _3062_ net941 _3747_ VGND VGND VPWR VPWR _3757_ sky130_fd_sc_hd__mux2_1
X_4814_ _1568_ _1569_ _1107_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__mux2_1
X_8582_ clknet_leaf_0_clk _0766_ VGND VGND VPWR VPWR rf.registers\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5794_ _2539_ _2540_ _2543_ VGND VGND VPWR VPWR _2544_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_32_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4644__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7533_ _3720_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4745_ _1499_ _1500_ _1259_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5745__A _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6340__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7464_ _3060_ net869 _3675_ VGND VGND VPWR VPWR _3684_ sky130_fd_sc_hd__mux2_1
X_4676_ rf.registers\[16\]\[22\] rf.registers\[17\]\[22\] rf.registers\[18\]\[22\]
+ rf.registers\[19\]\[22\] net135 _1184_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__mux4_1
XANTENNA__8160__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6415_ _3098_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9203_ clknet_leaf_34_clk _0363_ VGND VGND VPWR VPWR rf.registers\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_7395_ _3647_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9134_ clknet_leaf_43_clk _0294_ VGND VGND VPWR VPWR rf.registers\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6346_ _3050_ net431 _3044_ VGND VGND VPWR VPWR _3051_ sky130_fd_sc_hd__mux2_1
XANTENNA__8267__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9065_ clknet_leaf_51_clk _0225_ VGND VGND VPWR VPWR rf.registers\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6277_ _2621_ _2995_ _3001_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__o21bai_4
XFILLER_0_110_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8016_ _3976_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__clkbuf_1
X_5228_ rf.registers\[28\]\[26\] rf.registers\[29\]\[26\] rf.registers\[30\]\[26\]
+ rf.registers\[31\]\[26\] _1881_ _1883_ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5159_ _1913_ _1914_ _1889_ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__mux2_1
XANTENNA__4580__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8918_ clknet_leaf_24_clk _0078_ VGND VGND VPWR VPWR rf.registers\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8849_ clknet_leaf_43_clk _0009_ VGND VGND VPWR VPWR rf.registers\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4635__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7346__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5655__A _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4399__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5060__S1 _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4476__B1 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4323__S0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7110__A net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4874__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8390__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4530_ _1282_ _1285_ _1071_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold306 rf.registers\[3\]\[19\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _1171_ _1188_ _1216_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold317 rf.registers\[6\]\[25\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 rf.registers\[8\]\[6\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold339 rf.registers\[16\]\[19\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _2621_ _2921_ _2928_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__o21bai_2
XANTENNA__4703__A1 _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7180_ _3532_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4392_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6131_ _2586_ _2797_ VGND VGND VPWR VPWR _2863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6062_ _2040_ _2796_ _2797_ _2421_ VGND VGND VPWR VPWR _2798_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1006 rf.registers\[4\]\[5\] VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1017 rf.registers\[20\]\[30\] VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlygate4sd3_1
X_5013_ rf.registers\[8\]\[21\] rf.registers\[9\]\[21\] rf.registers\[10\]\[21\] rf.registers\[11\]\[21\]
+ _1767_ _1768_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__mux4_1
Xhold1028 rf.registers\[31\]\[19\] VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 rf.registers\[31\]\[9\] VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4562__S0 _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
X_6964_ _3402_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8703_ clknet_leaf_70_clk _0887_ VGND VGND VPWR VPWR rf.registers\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_5915_ _1464_ _2536_ _2658_ VGND VGND VPWR VPWR _2659_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6895_ net516 _3141_ _3362_ VGND VGND VPWR VPWR _3366_ sky130_fd_sc_hd__mux2_1
XANTENNA__8550__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5846_ _1060_ _1083_ VGND VGND VPWR VPWR _2594_ sky130_fd_sc_hd__nand2_1
X_8634_ clknet_leaf_37_clk _0818_ VGND VGND VPWR VPWR rf.registers\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8831__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6392__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5777_ _2524_ _2527_ _2501_ VGND VGND VPWR VPWR _2528_ sky130_fd_sc_hd__mux2_1
X_8565_ _4266_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7166__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5290__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7516_ _3043_ net639 _3711_ VGND VGND VPWR VPWR _3712_ sky130_fd_sc_hd__mux2_1
X_4728_ rf.registers\[20\]\[14\] rf.registers\[21\]\[14\] rf.registers\[22\]\[14\]
+ rf.registers\[23\]\[14\] _1324_ _1325_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__mux4_1
X_8496_ net477 net29 _4227_ VGND VGND VPWR VPWR _4231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7447_ _3663_ VGND VGND VPWR VPWR _3675_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4659_ _1025_ _1406_ _1410_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8981__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7378_ _3638_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
Xhold840 rf.registers\[13\]\[28\] VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold851 rf.registers\[30\]\[13\] VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold862 rf.registers\[1\]\[19\] VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 rf.registers\[12\]\[20\] VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__dlygate4sd3_1
X_6329_ net44 VGND VGND VPWR VPWR _3039_ sky130_fd_sc_hd__clkbuf_2
Xhold884 rf.registers\[31\]\[11\] VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__dlygate4sd3_1
X_9117_ clknet_leaf_3_clk _0277_ VGND VGND VPWR VPWR rf.registers\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold895 rf.registers\[21\]\[26\] VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__dlygate4sd3_1
X_9048_ clknet_leaf_12_clk _0208_ VGND VGND VPWR VPWR rf.registers\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7947__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4554__A _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4856__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8460__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8372__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6383__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5186__A1 _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5725__A3 _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5385__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7804__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6686__A1 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_max_cap81_A _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4544__S0 _1262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4464__A _1219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4847__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5700_ _2452_ _2453_ _2421_ VGND VGND VPWR VPWR _2454_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8370__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6680_ _3251_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5631_ _1167_ _2016_ VGND VGND VPWR VPWR _2386_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5295__A _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8350_ _4153_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__clkbuf_1
X_5562_ _1716_ _2317_ VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7301_ _3597_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4513_ rf.registers\[8\]\[21\] rf.registers\[9\]\[21\] rf.registers\[10\]\[21\] rf.registers\[11\]\[21\]
+ net1164 _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__mux4_1
X_8281_ _3130_ net726 _4108_ VGND VGND VPWR VPWR _4117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5493_ _1669_ _2230_ _2248_ VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__o21ai_1
Xhold103 rf.registers\[5\]\[25\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 rf.registers\[18\]\[16\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7232_ _3033_ net552 _3555_ VGND VGND VPWR VPWR _3561_ sky130_fd_sc_hd__mux2_1
Xhold125 rf.registers\[14\]\[10\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7874__A0 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4444_ _1027_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_7_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold136 rf.registers\[30\]\[12\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold147 rf.registers\[25\]\[26\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold158 rf.registers\[5\]\[8\] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold169 rf.registers\[20\]\[31\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ _3523_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
X_4375_ _1129_ _1130_ _1035_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__mux2_1
XANTENNA__4783__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5234__S _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6429__A1 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6114_ _2800_ _2847_ _1877_ VGND VGND VPWR VPWR _2848_ sky130_fd_sc_hd__mux2_1
X_7094_ _3480_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _1512_ _1602_ _1634_ _2658_ _2536_ VGND VGND VPWR VPWR _2782_ sky130_fd_sc_hd__a41o_1
XANTENNA__5101__A1 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ _3118_ net461 _3963_ VGND VGND VPWR VPWR _3966_ sky130_fd_sc_hd__mux2_1
XANTENNA__4838__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6947_ _3393_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6878_ net265 _3124_ _3351_ VGND VGND VPWR VPWR _3357_ sky130_fd_sc_hd__mux2_1
XANTENNA__8354__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8617_ clknet_leaf_51_clk _0801_ VGND VGND VPWR VPWR rf.registers\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5829_ _2418_ VGND VGND VPWR VPWR _2577_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5263__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4313__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8548_ net598 net21 _4255_ VGND VGND VPWR VPWR _4258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8479_ net792 net20 _4216_ VGND VGND VPWR VPWR _4222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4774__S0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold670 rf.registers\[28\]\[29\] VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5340__B2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold681 rf.registers\[16\]\[7\] VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold692 rf.registers\[12\]\[25\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7093__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4659__A1_N _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5643__A2 _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4284__A _1034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8190__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8345__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6004__A _1874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7534__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7856__A0 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5843__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5006__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output80_A net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4459__A _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5054__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5619__C1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4517__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4893__S _1645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6831__A1 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5190__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7850_ _3888_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__clkbuf_1
X_6801_ _3316_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6595__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7781_ net569 _3470_ _3844_ VGND VGND VPWR VPWR _3852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4993_ _1745_ _1746_ _1748_ _1697_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__o211a_1
XANTENNA__7709__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9520_ clknet_leaf_9_clk _0680_ VGND VGND VPWR VPWR rf.registers\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4922__A _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6732_ _3279_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6613__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6663_ net273 _3113_ _3242_ VGND VGND VPWR VPWR _3243_ sky130_fd_sc_hd__mux2_1
X_9451_ clknet_leaf_4_clk _0611_ VGND VGND VPWR VPWR rf.registers\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload69_A clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5245__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5614_ _1799_ _2306_ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__or2_1
X_8402_ _4181_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9382_ clknet_leaf_0_clk _0542_ VGND VGND VPWR VPWR rf.registers\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6594_ _3194_ VGND VGND VPWR VPWR _3206_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5545_ rf.registers\[4\]\[4\] rf.registers\[5\]\[4\] rf.registers\[6\]\[4\] rf.registers\[7\]\[4\]
+ _1718_ _1679_ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__mux4_1
X_8333_ net994 _3476_ _4144_ VGND VGND VPWR VPWR _4145_ sky130_fd_sc_hd__mux2_1
XANTENNA__7847__A0 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8264_ _4096_ VGND VGND VPWR VPWR _4108_ sky130_fd_sc_hd__buf_4
X_5476_ rf.registers\[28\]\[9\] rf.registers\[29\]\[9\] rf.registers\[30\]\[9\] rf.registers\[31\]\[9\]
+ _1675_ _1692_ VGND VGND VPWR VPWR _2232_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4427_ _1044_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__buf_4
X_7215_ _3550_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_8195_ _4071_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7146_ net309 _3450_ _3455_ VGND VGND VPWR VPWR _3514_ sky130_fd_sc_hd__mux2_1
X_4358_ rf.registers\[16\]\[2\] rf.registers\[17\]\[2\] rf.registers\[18\]\[2\] rf.registers\[19\]\[2\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_6_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ net913 _3468_ _3456_ VGND VGND VPWR VPWR _3469_ sky130_fd_sc_hd__mux2_1
XANTENNA__8275__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4508__S0 _1262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4289_ rf.registers\[4\]\[4\] rf.registers\[5\]\[4\] rf.registers\[6\]\[4\] rf.registers\[7\]\[4\]
+ net103 _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__mux4_1
X_6028_ _2755_ _2760_ _2766_ _2621_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_87_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4308__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7979_ _3101_ net741 _3952_ VGND VGND VPWR VPWR _3957_ sky130_fd_sc_hd__mux2_1
XANTENNA__7619__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6889__A1 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4995__S0 _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7354__S _3590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4279__A _1034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4747__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5172__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8015__A0 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4521__A1_N _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8566__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5475__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload12 clknet_leaf_71_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_153_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload23 clknet_leaf_65_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__4986__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload34 clknet_leaf_46_clk VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__inv_8
XANTENNA__7264__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload45 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__inv_6
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5330_ rf.registers\[16\]\[1\] rf.registers\[17\]\[1\] rf.registers\[18\]\[1\] rf.registers\[19\]\[1\]
+ _1673_ _1690_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload56 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload56/Y sky130_fd_sc_hd__clkinv_8
Xclkload67 clknet_leaf_31_clk VGND VGND VPWR VPWR clkload67/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_53_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5261_ _1668_ _2016_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_149_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7000_ net236 _3109_ _3413_ VGND VGND VPWR VPWR _3422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5192_ rf.registers\[20\]\[28\] rf.registers\[21\]\[28\] rf.registers\[22\]\[28\]
+ rf.registers\[23\]\[28\] _1882_ _1884_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_118_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8254__A0 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4917__A _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8951_ clknet_leaf_23_clk _0111_ VGND VGND VPWR VPWR rf.registers\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4815__B1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7902_ _3915_ VGND VGND VPWR VPWR _3916_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8882_ clknet_leaf_37_clk _0042_ VGND VGND VPWR VPWR rf.registers\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7833_ _3021_ _3193_ VGND VGND VPWR VPWR _3879_ sky130_fd_sc_hd__nand2_4
XFILLER_0_66_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7439__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5466__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6343__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7764_ _3842_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_82_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4976_ _1639_ _1731_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_127_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9503_ clknet_leaf_71_clk _0663_ VGND VGND VPWR VPWR rf.registers\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6715_ _3270_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4371__B _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7695_ net831 _3452_ _3771_ VGND VGND VPWR VPWR _3806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5218__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9434_ clknet_leaf_17_clk _0594_ VGND VGND VPWR VPWR rf.registers\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xclkload6 clknet_3_7__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinvlp_4
X_6646_ net1048 _3097_ _3231_ VGND VGND VPWR VPWR _3234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9365_ clknet_leaf_35_clk _0525_ VGND VGND VPWR VPWR rf.registers\[20\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6577_ _3197_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8316_ net835 _3460_ _4133_ VGND VGND VPWR VPWR _4136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5528_ _2282_ _2283_ _1738_ VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__mux2_1
X_9296_ clknet_leaf_4_clk _0456_ VGND VGND VPWR VPWR rf.registers\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ rf.registers\[16\]\[8\] rf.registers\[17\]\[8\] rf.registers\[18\]\[8\] rf.registers\[19\]\[8\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2215_ sky130_fd_sc_hd__mux4_1
X_8247_ _4099_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4729__S0 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8178_ net150 _3458_ _4061_ VGND VGND VPWR VPWR _4063_ sky130_fd_sc_hd__mux2_1
XANTENNA__7048__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6518__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7129_ net29 VGND VGND VPWR VPWR _3504_ sky130_fd_sc_hd__buf_2
XANTENNA__5154__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4901__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8548__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5782__A1 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6731__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4968__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5393__S0 _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7113__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8539__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8595__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7259__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5568__A _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4830_ _1205_ _1585_ _1170_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ rf.registers\[24\]\[8\] rf.registers\[25\]\[8\] rf.registers\[26\]\[8\] rf.registers\[27\]\[8\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6500_ net10 net9 net46 VGND VGND VPWR VPWR _3154_ sky130_fd_sc_hd__or3b_1
X_7480_ _3692_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
X_4692_ net122 _1447_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6431_ net44 VGND VGND VPWR VPWR _3109_ sky130_fd_sc_hd__buf_2
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9150_ clknet_leaf_0_clk _0310_ VGND VGND VPWR VPWR rf.registers\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6362_ _3061_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__clkbuf_1
X_5313_ rf.registers\[24\]\[2\] rf.registers\[25\]\[2\] rf.registers\[26\]\[2\] rf.registers\[27\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2069_ sky130_fd_sc_hd__mux4_1
X_8101_ _4021_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6293_ net301 _3013_ _3007_ VGND VGND VPWR VPWR _3014_ sky130_fd_sc_hd__mux2_1
X_9081_ clknet_leaf_19_clk _0241_ VGND VGND VPWR VPWR rf.registers\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7722__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8032_ _3984_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__clkbuf_1
X_5244_ rf.registers\[20\]\[25\] rf.registers\[21\]\[25\] rf.registers\[22\]\[25\]
+ rf.registers\[23\]\[25\] _1822_ _1823_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__mux4_1
XANTENNA__4500__A2 _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5175_ rf.registers\[24\]\[29\] rf.registers\[25\]\[29\] rf.registers\[26\]\[29\]
+ rf.registers\[27\]\[29\] _1705_ _1708_ VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__mux4_1
XANTENNA__5136__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8934_ clknet_leaf_2_clk _0094_ VGND VGND VPWR VPWR rf.registers\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8865_ clknet_leaf_56_clk _0025_ VGND VGND VPWR VPWR rf.registers\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5439__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7816_ _3870_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8796_ clknet_leaf_16_clk _0980_ VGND VGND VPWR VPWR rf.registers\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7747_ _3071_ net538 _3830_ VGND VGND VPWR VPWR _3834_ sky130_fd_sc_hd__mux2_1
X_4959_ _1700_ _1714_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7678_ _3797_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_1
X_9417_ clknet_leaf_45_clk _0577_ VGND VGND VPWR VPWR rf.registers\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6629_ _3224_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5417__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9348_ clknet_leaf_52_clk _0508_ VGND VGND VPWR VPWR rf.registers\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_95_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9279_ clknet_leaf_73_clk _0439_ VGND VGND VPWR VPWR rf.registers\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6248__S _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5152__S _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4350__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5388__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4292__A _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5062__S _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4494__A1 _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6980_ _3410_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5931_ _1800_ _2194_ _2176_ VGND VGND VPWR VPWR _2675_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5994__A1 _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8650_ clknet_leaf_7_clk _0834_ VGND VGND VPWR VPWR rf.registers\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_5862_ _2353_ _2358_ VGND VGND VPWR VPWR _2609_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7601_ _3756_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4813_ rf.registers\[0\]\[11\] rf.registers\[1\]\[11\] rf.registers\[2\]\[11\] rf.registers\[3\]\[11\]
+ net102 _1090_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__mux4_1
X_8581_ clknet_leaf_62_clk _0765_ VGND VGND VPWR VPWR rf.registers\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5793_ _2511_ _2512_ _2518_ _2542_ VGND VGND VPWR VPWR _2543_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_56_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7717__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4930__A _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7532_ _3060_ net425 _3711_ VGND VGND VPWR VPWR _3720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4744_ rf.registers\[24\]\[15\] rf.registers\[25\]\[15\] rf.registers\[26\]\[15\]
+ rf.registers\[27\]\[15\] _1324_ _1325_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__mux4_1
XANTENNA__5745__B _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7463_ _3683_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_1
X_4675_ rf.registers\[20\]\[22\] rf.registers\[21\]\[22\] rf.registers\[22\]\[22\]
+ rf.registers\[23\]\[22\] net135 _1184_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9202_ clknet_leaf_42_clk _0362_ VGND VGND VPWR VPWR rf.registers\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6414_ net436 _3097_ _3093_ VGND VGND VPWR VPWR _3098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7394_ _3058_ net880 _3639_ VGND VGND VPWR VPWR _3647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9133_ clknet_leaf_50_clk _0293_ VGND VGND VPWR VPWR rf.registers\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6345_ net18 VGND VGND VPWR VPWR _3050_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__8548__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7452__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9064_ clknet_leaf_49_clk _0224_ VGND VGND VPWR VPWR rf.registers\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6276_ _2720_ _2737_ _2996_ _2472_ _3000_ VGND VGND VPWR VPWR _3001_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5227_ _1981_ _1982_ _1901_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__mux2_1
X_8015_ _3137_ net773 _3974_ VGND VGND VPWR VPWR _3976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5109__S0 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5158_ rf.registers\[12\]\[30\] rf.registers\[13\]\[30\] rf.registers\[14\]\[30\]
+ rf.registers\[15\]\[30\] _1881_ _1883_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__mux4_1
XANTENNA__4580__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8283__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5089_ _1843_ _1844_ _1686_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8917_ clknet_leaf_32_clk _0077_ VGND VGND VPWR VPWR rf.registers\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8848_ clknet_leaf_10_clk _0008_ VGND VGND VPWR VPWR rf.registers\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8779_ clknet_leaf_4_clk _0963_ VGND VGND VPWR VPWR rf.registers\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7627__S _3735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6531__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4840__A _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4399__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8458__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7662__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4476__A1 _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6706__S _3230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4323__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5520__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5846__A _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7537__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4750__A _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4460_ _1197_ _1206_ _1212_ _1214_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__o221a_4
XTAP_TAPCELL_ROW_152_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold307 rf.registers\[13\]\[30\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7350__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold318 rf.registers\[7\]\[2\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold329 rf.registers\[3\]\[2\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5082__A1_N _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8368__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4391_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__7272__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5581__A _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6130_ _2621_ _2856_ _2862_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__o21a_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4909__B _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6061_ _2737_ VGND VGND VPWR VPWR _2797_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9139__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _1707_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__clkbuf_4
Xhold1007 rf.registers\[4\]\[23\] VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 rf.registers\[24\]\[22\] VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 rf.registers\[20\]\[21\] VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6616__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4925__A _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5511__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6963_ net1089 _3141_ _3398_ VGND VGND VPWR VPWR _3402_ sky130_fd_sc_hd__mux2_1
X_8702_ clknet_leaf_71_clk _0886_ VGND VGND VPWR VPWR rf.registers\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_5914_ _2657_ VGND VGND VPWR VPWR _2658_ sky130_fd_sc_hd__buf_6
XFILLER_0_76_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6894_ _3365_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8633_ clknet_leaf_20_clk _0817_ VGND VGND VPWR VPWR rf.registers\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5845_ _1111_ net83 _1145_ net1168 VGND VGND VPWR VPWR _2593_ sky130_fd_sc_hd__nand4_2
XFILLER_0_146_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5756__A _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8564_ net1137 net30 _3006_ VGND VGND VPWR VPWR _4266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ _2363_ _2456_ _2526_ VGND VGND VPWR VPWR _2527_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7515_ _3699_ VGND VGND VPWR VPWR _3711_ sky130_fd_sc_hd__buf_4
X_4727_ rf.registers\[16\]\[14\] rf.registers\[17\]\[14\] rf.registers\[18\]\[14\]
+ rf.registers\[19\]\[14\] _1324_ _1325_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8495_ _4230_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7446_ _3674_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__clkbuf_1
X_4658_ _1078_ _1413_ _1057_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold830 rf.registers\[29\]\[29\] VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__dlygate4sd3_1
X_7377_ _3041_ net1085 _3628_ VGND VGND VPWR VPWR _3638_ sky130_fd_sc_hd__mux2_1
Xhold841 rf.registers\[8\]\[24\] VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5491__A _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold852 rf.registers\[15\]\[16\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd3_1
X_4589_ rf.registers\[0\]\[30\] rf.registers\[1\]\[30\] rf.registers\[2\]\[30\] rf.registers\[3\]\[30\]
+ net128 _1263_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9116_ clknet_leaf_16_clk _0276_ VGND VGND VPWR VPWR rf.registers\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold863 rf.registers\[30\]\[28\] VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 rf.registers\[16\]\[25\] VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ _3038_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__clkbuf_1
Xhold885 rf.registers\[23\]\[28\] VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 rf.registers\[18\]\[22\] VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9047_ clknet_leaf_33_clk _0207_ VGND VGND VPWR VPWR rf.registers\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6259_ _1923_ _2983_ VGND VGND VPWR VPWR _2985_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_123_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5958__A1 _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clone35_A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7332__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8188__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4544__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8217__A _4060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5576__A _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5630_ _2383_ _2384_ VGND VGND VPWR VPWR _2385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5561_ _2315_ _2316_ _1711_ VGND VGND VPWR VPWR _2317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7300_ _3033_ net1007 _3591_ VGND VGND VPWR VPWR _3597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7323__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4512_ _1202_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__buf_4
X_5492_ _1668_ _2247_ VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__nand2_1
X_8280_ _4116_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold104 rf.registers\[10\]\[27\] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 rf.registers\[6\]\[8\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7231_ _3560_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
Xhold126 rf.registers\[7\]\[17\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4443_ _1198_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__buf_4
XANTENNA__8098__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold137 rf.registers\[8\]\[0\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 rf.registers\[11\]\[13\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5885__B1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold159 rf.registers\[3\]\[27\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
X_7162_ net282 _3466_ _3517_ VGND VGND VPWR VPWR _3523_ sky130_fd_sc_hd__mux2_1
X_4374_ rf.registers\[16\]\[1\] rf.registers\[17\]\[1\] rf.registers\[18\]\[1\] rf.registers\[19\]\[1\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux4_2
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4783__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6113_ _1781_ _1756_ VGND VGND VPWR VPWR _2847_ sky130_fd_sc_hd__and2_1
X_7093_ net943 _3479_ _3477_ VGND VGND VPWR VPWR _3480_ sky130_fd_sc_hd__mux2_1
XANTENNA__7730__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6044_ _2408_ _2775_ _2776_ _2781_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__o22a_1
XANTENNA__6346__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5250__S _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7995_ _3965_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4299__S0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6062__B1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6946_ net535 _3124_ _3387_ VGND VGND VPWR VPWR _3393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6877_ _3356_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7177__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5486__A _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8616_ clknet_leaf_52_clk _0800_ VGND VGND VPWR VPWR rf.registers\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4390__A _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5828_ _2504_ _2564_ _2576_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__a21o_1
XFILLER_0_64_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8547_ _4257_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__clkbuf_1
X_5759_ _2509_ _2510_ VGND VGND VPWR VPWR _2511_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7905__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8478_ _4221_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7429_ _3025_ net1124 _3664_ VGND VGND VPWR VPWR _3666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold660 rf.registers\[31\]\[28\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 rf.registers\[2\]\[9\] VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4774__S1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold682 rf.registers\[10\]\[7\] VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold693 rf.registers\[16\]\[21\] VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7876__A _3879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8471__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4504__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7553__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4462__S0 _1182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7815__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5843__B _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7116__A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6020__A _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output73_A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4517__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5190__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6800_ net177 _3113_ _3315_ VGND VGND VPWR VPWR _3316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7780_ _3851_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__clkbuf_1
X_4992_ _1712_ _1747_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6731_ _3043_ net207 _3278_ VGND VGND VPWR VPWR _3279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9450_ clknet_leaf_7_clk _0610_ VGND VGND VPWR VPWR rf.registers\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6662_ _3230_ VGND VGND VPWR VPWR _3242_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8401_ net286 _3476_ _4180_ VGND VGND VPWR VPWR _4181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_5613_ _1167_ _2063_ VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__nand2_1
X_9381_ clknet_leaf_57_clk _0541_ VGND VGND VPWR VPWR rf.registers\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6593_ _3205_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4453__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8332_ _4132_ VGND VGND VPWR VPWR _4144_ sky130_fd_sc_hd__clkbuf_8
X_5544_ _1716_ _2299_ VGND VGND VPWR VPWR _2300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8263_ _4107_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5475_ rf.registers\[24\]\[9\] rf.registers\[25\]\[9\] rf.registers\[26\]\[9\] rf.registers\[27\]\[9\]
+ _1675_ _1692_ VGND VGND VPWR VPWR _2231_ sky130_fd_sc_hd__mux4_1
X_7214_ net287 _3450_ _3516_ VGND VGND VPWR VPWR _3550_ sky130_fd_sc_hd__mux2_1
X_4426_ net1155 VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__buf_12
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8194_ net143 _3474_ _4061_ VGND VGND VPWR VPWR _4071_ sky130_fd_sc_hd__mux2_1
XANTENNA__8556__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7145_ _3513_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
X_4357_ rf.registers\[28\]\[2\] rf.registers\[29\]\[2\] rf.registers\[30\]\[2\] rf.registers\[31\]\[2\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_6_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7460__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7076_ net42 VGND VGND VPWR VPWR _3468_ sky130_fd_sc_hd__buf_2
X_4288_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__buf_4
XANTENNA__4508__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6027_ _2763_ _2765_ VGND VGND VPWR VPWR _2766_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_87_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6804__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7978_ _3956_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ net974 _3107_ _3376_ VGND VGND VPWR VPWR _3384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6105__A _1754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9579_ clknet_leaf_5_clk _0739_ VGND VGND VPWR VPWR rf.registers\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7635__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4995__S1 _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5155__S _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6510__A1 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4747__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold490 rf.registers\[15\]\[13\] VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8466__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5172__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6714__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7526__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5001__A1 _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7545__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload13 clknet_leaf_72_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_6
XFILLER_0_113_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload24 clknet_leaf_52_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_152_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload35 clknet_leaf_47_clk VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__inv_6
XANTENNA__4986__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload46 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload46/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_2_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload57 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload57/Y sky130_fd_sc_hd__clkinv_8
Xclkload68 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload68/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5260_ net1163 _2015_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8376__S _4132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5191_ rf.registers\[16\]\[28\] rf.registers\[17\]\[28\] rf.registers\[18\]\[28\]
+ rf.registers\[19\]\[28\] _1882_ _1884_ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__mux4_1
XANTENNA__7280__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6265__B1 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8950_ clknet_leaf_24_clk _0110_ VGND VGND VPWR VPWR rf.registers\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4815__A1 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7901_ _3005_ _3090_ VGND VGND VPWR VPWR _3915_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_69_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8881_ clknet_leaf_39_clk _0041_ VGND VGND VPWR VPWR rf.registers\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6624__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7832_ _3878_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4933__A _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7763_ _3087_ net603 _3807_ VGND VGND VPWR VPWR _3842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4975_ _1672_ _1698_ _1715_ _1730_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_82_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5240__A1 _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9502_ clknet_leaf_71_clk _0662_ VGND VGND VPWR VPWR rf.registers\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6714_ _3027_ net857 _3267_ VGND VGND VPWR VPWR _3270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7694_ _3805_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9433_ clknet_leaf_20_clk _0593_ VGND VGND VPWR VPWR rf.registers\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6645_ _3233_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__clkbuf_1
Xclkload7 clknet_leaf_66_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9364_ clknet_leaf_38_clk _0524_ VGND VGND VPWR VPWR rf.registers\[20\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6576_ _3025_ net970 _3195_ VGND VGND VPWR VPWR _3197_ sky130_fd_sc_hd__mux2_1
XANTENNA__8867__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8315_ _4135_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__clkbuf_1
X_5527_ rf.registers\[0\]\[7\] rf.registers\[1\]\[7\] rf.registers\[2\]\[7\] rf.registers\[3\]\[7\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9295_ clknet_leaf_9_clk _0455_ VGND VGND VPWR VPWR rf.registers\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8246_ _3095_ net707 _4097_ VGND VGND VPWR VPWR _4099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5458_ rf.registers\[20\]\[8\] rf.registers\[21\]\[8\] rf.registers\[22\]\[8\] rf.registers\[23\]\[8\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2214_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4729__S1 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4409_ _1088_ _1164_ net8 VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a21oi_2
XANTENNA__8286__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8177_ _4062_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__clkbuf_1
X_5389_ rf.registers\[20\]\[13\] rf.registers\[21\]\[13\] rf.registers\[22\]\[13\]
+ rf.registers\[23\]\[13\] _1673_ _1690_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7128_ _3503_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7059_ net506 _3454_ _3456_ VGND VGND VPWR VPWR _3457_ sky130_fd_sc_hd__mux2_1
XANTENNA__5154__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4901__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4665__S0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_rebuffer45_A _1166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7365__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5674__A _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4968__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5090__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5393__S1 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8236__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5568__B _2323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4656__S0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ rf.registers\[28\]\[8\] rf.registers\[29\]\[8\] rf.registers\[30\]\[8\] rf.registers\[31\]\[8\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_16_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4691_ _1430_ _1446_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__and2_4
XFILLER_0_153_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6430_ _3108_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4733__B1 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6361_ _3060_ net433 _3044_ VGND VGND VPWR VPWR _3061_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8100_ net965 _3448_ _4011_ VGND VGND VPWR VPWR _4021_ sky130_fd_sc_hd__mux2_1
X_5312_ rf.registers\[28\]\[2\] rf.registers\[29\]\[2\] rf.registers\[30\]\[2\] rf.registers\[31\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__mux4_1
XANTENNA__8475__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9080_ clknet_leaf_11_clk _0240_ VGND VGND VPWR VPWR rf.registers\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6292_ net35 VGND VGND VPWR VPWR _3013_ sky130_fd_sc_hd__clkbuf_4
X_8031_ _3013_ net1118 _3974_ VGND VGND VPWR VPWR _3984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5243_ _1980_ _1998_ VGND VGND VPWR VPWR _1999_ sky130_fd_sc_hd__or2_1
XANTENNA__4928__A _1645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5174_ rf.registers\[28\]\[29\] rf.registers\[29\]\[29\] rf.registers\[30\]\[29\]
+ rf.registers\[31\]\[29\] _1705_ _1708_ VGND VGND VPWR VPWR _1930_ sky130_fd_sc_hd__mux4_1
XANTENNA__6789__A1 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5136__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8933_ clknet_leaf_52_clk _0093_ VGND VGND VPWR VPWR rf.registers\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4895__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8864_ clknet_leaf_69_clk _0024_ VGND VGND VPWR VPWR rf.registers\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7738__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7815_ net153 _3504_ _3866_ VGND VGND VPWR VPWR _3870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8795_ clknet_leaf_22_clk _0979_ VGND VGND VPWR VPWR rf.registers\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4647__S0 _1104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7746_ _3833_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4958_ _1709_ _1710_ _1713_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7677_ net582 _3502_ _3794_ VGND VGND VPWR VPWR _3797_ sky130_fd_sc_hd__mux2_1
X_4889_ net3 VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__inv_2
XANTENNA__7185__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4602__S _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9416_ clknet_leaf_45_clk _0576_ VGND VGND VPWR VPWR rf.registers\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6628_ _3077_ net492 _3217_ VGND VGND VPWR VPWR _3224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9347_ clknet_leaf_61_clk _0507_ VGND VGND VPWR VPWR rf.registers\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6559_ _3186_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7913__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8466__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9278_ clknet_leaf_73_clk _0438_ VGND VGND VPWR VPWR rf.registers\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8229_ _4089_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6529__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8218__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7977__A0 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_67_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7823__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6439__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8209__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5930_ _2212_ _2429_ VGND VGND VPWR VPWR _2674_ sky130_fd_sc_hd__nor2_1
XANTENNA__4483__A _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5861_ _2457_ _2525_ _1877_ VGND VGND VPWR VPWR _2608_ sky130_fd_sc_hd__mux2_1
XANTENNA__7196__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7600_ _3060_ net801 _3747_ VGND VGND VPWR VPWR _3756_ sky130_fd_sc_hd__mux2_1
X_4812_ rf.registers\[4\]\[11\] rf.registers\[5\]\[11\] rf.registers\[6\]\[11\] rf.registers\[7\]\[11\]
+ net102 _1090_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__mux4_1
X_8580_ clknet_leaf_62_clk _0764_ VGND VGND VPWR VPWR rf.registers\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5792_ _2509_ _2541_ _2517_ VGND VGND VPWR VPWR _2542_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7531_ _3719_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4743_ rf.registers\[28\]\[15\] rf.registers\[29\]\[15\] rf.registers\[30\]\[15\]
+ rf.registers\[31\]\[15\] net128 _1263_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7462_ _3058_ net972 _3675_ VGND VGND VPWR VPWR _3683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4674_ _1239_ _1421_ _1425_ _1429_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__a2bb2o_2
X_9201_ clknet_leaf_40_clk _0361_ VGND VGND VPWR VPWR rf.registers\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6413_ net36 VGND VGND VPWR VPWR _3097_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7393_ _3646_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9132_ clknet_leaf_50_clk _0292_ VGND VGND VPWR VPWR rf.registers\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8448__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6344_ _3049_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9063_ clknet_leaf_65_clk _0223_ VGND VGND VPWR VPWR rf.registers\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6349__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6275_ _2530_ _2859_ _2999_ _1087_ VGND VGND VPWR VPWR _3000_ sky130_fd_sc_hd__o211a_1
XANTENNA__5253__S _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8014_ _3975_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__clkbuf_1
X_5226_ rf.registers\[16\]\[26\] rf.registers\[17\]\[26\] rf.registers\[18\]\[26\]
+ rf.registers\[19\]\[26\] _1881_ _1883_ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_90_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5682__A1 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8564__S _3006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5157_ rf.registers\[8\]\[30\] rf.registers\[9\]\[30\] rf.registers\[10\]\[30\] rf.registers\[11\]\[30\]
+ _1881_ _1883_ VGND VGND VPWR VPWR _1913_ sky130_fd_sc_hd__mux4_1
XANTENNA__5109__S1 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5088_ rf.registers\[16\]\[17\] rf.registers\[17\]\[17\] rf.registers\[18\]\[17\]
+ rf.registers\[19\]\[17\] _1689_ _1693_ VGND VGND VPWR VPWR _1844_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_108_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8916_ clknet_leaf_29_clk _0076_ VGND VGND VPWR VPWR rf.registers\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4642__C1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8847_ clknet_leaf_29_clk _0007_ VGND VGND VPWR VPWR rf.registers\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6812__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8778_ clknet_leaf_7_clk _0962_ VGND VGND VPWR VPWR rf.registers\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7729_ _3824_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7643__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5952__A _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4568__A _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4859__S0 _1173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5520__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__9210__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6722__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6925__A1 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_154_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7119__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6023__A _1601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5036__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold308 rf.registers\[21\]\[15\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7553__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold319 rf.registers\[18\]\[8\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4390_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_59_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5581__B _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7102__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6060_ _2585_ _2578_ _2426_ VGND VGND VPWR VPWR _2796_ sky130_fd_sc_hd__mux2_1
Xhold1008 rf.registers\[25\]\[11\] VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _1704_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__buf_4
XANTENNA__8384__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 rf.registers\[21\]\[1\] VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6613__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6962_ _3401_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5967__A2 _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5511__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5913_ _1416_ _1573_ _2506_ _2535_ VGND VGND VPWR VPWR _2657_ sky130_fd_sc_hd__and4b_2
X_8701_ clknet_leaf_15_clk _0885_ VGND VGND VPWR VPWR rf.registers\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6893_ net403 _3139_ _3362_ VGND VGND VPWR VPWR _3365_ sky130_fd_sc_hd__mux2_1
XANTENNA__7728__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6632__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8632_ clknet_leaf_27_clk _0816_ VGND VGND VPWR VPWR rf.registers\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4941__A _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5844_ _2038_ _2590_ _2591_ _2253_ VGND VGND VPWR VPWR _2592_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_118_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8563_ _4265_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__clkbuf_1
X_5775_ _2327_ _2525_ VGND VGND VPWR VPWR _2526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7514_ _3710_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_79_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4726_ rf.registers\[28\]\[14\] rf.registers\[29\]\[14\] rf.registers\[30\]\[14\]
+ rf.registers\[31\]\[14\] _1324_ _1325_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__mux4_1
XANTENNA__6129__C1 _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8494_ net647 net28 _4227_ VGND VGND VPWR VPWR _4230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5027__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7445_ _3041_ net954 _3664_ VGND VGND VPWR VPWR _3674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4657_ _1411_ _1412_ _1040_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold820 rf.registers\[16\]\[29\] VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd3_1
X_7376_ _3637_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_92_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold831 rf.registers\[3\]\[6\] VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4588_ rf.registers\[4\]\[30\] rf.registers\[5\]\[30\] rf.registers\[6\]\[30\] rf.registers\[7\]\[30\]
+ net128 _1263_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__mux4_1
Xhold842 rf.registers\[2\]\[0\] VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5491__B _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold853 rf.registers\[15\]\[10\] VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd3_1
X_9115_ clknet_leaf_36_clk _0275_ VGND VGND VPWR VPWR rf.registers\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6327_ _3037_ net905 _3023_ VGND VGND VPWR VPWR _3038_ sky130_fd_sc_hd__mux2_1
Xhold864 rf.registers\[12\]\[15\] VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold875 rf.registers\[30\]\[14\] VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold886 rf.registers\[3\]\[15\] VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 rf.registers\[27\]\[23\] VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__dlygate4sd3_1
X_9046_ clknet_leaf_24_clk _0206_ VGND VGND VPWR VPWR rf.registers\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6258_ _1923_ _2983_ VGND VGND VPWR VPWR _2984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8294__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5209_ _1963_ _1964_ _1745_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__mux2_1
X_6189_ _2916_ _2917_ VGND VGND VPWR VPWR _2918_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5012__A _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6907__A1 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5266__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5772__A1_N _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5018__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8469__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6778__A _3303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7373__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkload0_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5857__A _2390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5576__B _1660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5560_ rf.registers\[12\]\[5\] rf.registers\[13\]\[5\] rf.registers\[14\]\[5\] rf.registers\[15\]\[5\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2316_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4511_ _1200_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__buf_12
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5491_ _1842_ _2246_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7230_ _3031_ net493 _3555_ VGND VGND VPWR VPWR _3560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold105 rf.registers\[10\]\[13\] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ _1040_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__buf_4
Xhold116 rf.registers\[9\]\[29\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 rf.registers\[0\]\[0\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 rf.registers\[3\]\[8\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold149 rf.registers\[0\]\[6\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7161_ _3522_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4373_ rf.registers\[20\]\[1\] rf.registers\[21\]\[1\] rf.registers\[22\]\[1\] rf.registers\[23\]\[1\]
+ net101 _1066_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__mux4_2
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6112_ _2102_ _2554_ VGND VGND VPWR VPWR _2846_ sky130_fd_sc_hd__nor2_1
X_7092_ net16 VGND VGND VPWR VPWR _3479_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6043_ _2625_ _2731_ _2779_ _2496_ _2780_ VGND VGND VPWR VPWR _2781_ sky130_fd_sc_hd__a221o_1
XANTENNA__4936__A _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7994_ _3116_ rf.registers\[21\]\[11\] _3963_ VGND VGND VPWR VPWR _3965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4299__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6062__A1 _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6945_ _3392_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7458__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6876_ net199 _3122_ _3351_ VGND VGND VPWR VPWR _3356_ sky130_fd_sc_hd__mux2_1
XANTENNA__5248__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8615_ clknet_leaf_63_clk _0799_ VGND VGND VPWR VPWR rf.registers\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5827_ _2496_ _2569_ _2572_ _2468_ _2575_ VGND VGND VPWR VPWR _2576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5758_ _2305_ _2508_ VGND VGND VPWR VPWR _2510_ sky130_fd_sc_hd__and2_1
XANTENNA__5573__B1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8546_ net472 net20 _4255_ VGND VGND VPWR VPWR _4257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4709_ rf.registers\[20\]\[13\] rf.registers\[21\]\[13\] rf.registers\[22\]\[13\]
+ rf.registers\[23\]\[13\] net126 _1029_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__mux4_1
X_8477_ net192 net19 _4216_ VGND VGND VPWR VPWR _4221_ sky130_fd_sc_hd__mux2_1
X_5689_ _1961_ _1999_ _2347_ VGND VGND VPWR VPWR _2443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7428_ _3665_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_116_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5876__A1 _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7359_ _3019_ net463 _3628_ VGND VGND VPWR VPWR _3629_ sky130_fd_sc_hd__mux2_1
Xhold650 rf.registers\[14\]\[20\] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 rf.registers\[12\]\[11\] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7921__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold672 rf.registers\[4\]\[14\] VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 rf.registers\[15\]\[21\] VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 rf.registers\[15\]\[24\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd3_1
X_9029_ clknet_leaf_61_clk _0189_ VGND VGND VPWR VPWR rf.registers\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6537__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5441__S _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6053__A1 _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5487__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone50 _1172_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_16
XANTENNA__4462__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8199__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6301__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5411__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7831__S _3843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5619__A1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output66_A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7132__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6044__A1 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5478__S0 _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4991_ rf.registers\[8\]\[22\] rf.registers\[9\]\[22\] rf.registers\[10\]\[22\] rf.registers\[11\]\[22\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__mux4_1
XANTENNA__7278__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5587__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6730_ _3266_ VGND VGND VPWR VPWR _3278_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ _3241_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5612_ _1167_ _2081_ VGND VGND VPWR VPWR _2367_ sky130_fd_sc_hd__or2_1
X_8400_ _4168_ VGND VGND VPWR VPWR _4180_ sky130_fd_sc_hd__buf_4
X_9380_ clknet_leaf_62_clk _0540_ VGND VGND VPWR VPWR rf.registers\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6592_ _3041_ net607 _3195_ VGND VGND VPWR VPWR _3205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4453__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8331_ _4143_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__clkbuf_1
X_5543_ _2297_ _2298_ _1738_ VGND VGND VPWR VPWR _2299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4430__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8262_ _3111_ net428 _4097_ VGND VGND VPWR VPWR _4107_ sky130_fd_sc_hd__mux2_1
X_5474_ _1639_ _2229_ VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__or2_1
X_7213_ _3549_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
X_4425_ _1042_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__buf_12
XFILLER_0_100_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8193_ _4070_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7741__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7144_ net430 _3448_ _3498_ VGND VGND VPWR VPWR _3513_ sky130_fd_sc_hd__mux2_1
X_4356_ rf.registers\[24\]\[2\] rf.registers\[25\]\[2\] rf.registers\[26\]\[2\] rf.registers\[27\]\[2\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__mux4_2
XFILLER_0_111_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _3467_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
X_4287_ A2[1] VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__buf_4
X_6026_ _2744_ _2749_ _2764_ VGND VGND VPWR VPWR _2765_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6035__A1 _1858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5469__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7977_ _3099_ net402 _3952_ VGND VGND VPWR VPWR _3956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ _3383_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6859_ net257 _3105_ _3340_ VGND VGND VPWR VPWR _3347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9578_ clknet_leaf_7_clk _0738_ VGND VGND VPWR VPWR rf.registers\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8529_ net764 net43 _4244_ VGND VGND VPWR VPWR _4248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6121__A _1731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__9571__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold480 rf.registers\[20\]\[16\] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 rf.registers\[20\]\[13\] VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6274__B2 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4380__S0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4515__S _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload14 clknet_leaf_73_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload25 clknet_leaf_53_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__inv_12
XFILLER_0_113_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload36 clknet_leaf_48_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__inv_12
XFILLER_0_152_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6031__A _1820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload47 clknet_leaf_14_clk VGND VGND VPWR VPWR clkload47/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload58 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload58/Y sky130_fd_sc_hd__inv_8
Xclkload69 clknet_leaf_35_clk VGND VGND VPWR VPWR clkload69/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5870__A _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5190_ rf.registers\[28\]\[28\] rf.registers\[29\]\[28\] rf.registers\[30\]\[28\]
+ rf.registers\[31\]\[28\] _1882_ _1884_ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__mux4_1
XANTENNA__8392__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7900_ _3914_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6905__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8880_ clknet_leaf_13_clk _0040_ VGND VGND VPWR VPWR rf.registers\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7831_ net168 _3452_ _3843_ VGND VGND VPWR VPWR _3878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7762_ _3841_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__clkbuf_1
X_4974_ _1717_ _1727_ _1729_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9501_ clknet_leaf_13_clk _0661_ VGND VGND VPWR VPWR rf.registers\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6713_ _3269_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__clkbuf_1
X_7693_ net736 _3450_ _3771_ VGND VGND VPWR VPWR _3805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7736__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6644_ net860 _3095_ _3231_ VGND VGND VPWR VPWR _3233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9432_ clknet_leaf_11_clk _0592_ VGND VGND VPWR VPWR rf.registers\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8421__A _4168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_67_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__8190__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6575_ _3196_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__clkbuf_1
X_9363_ clknet_leaf_36_clk _0523_ VGND VGND VPWR VPWR rf.registers\[20\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8314_ net405 _3458_ _4133_ VGND VGND VPWR VPWR _4135_ sky130_fd_sc_hd__mux2_1
X_5526_ rf.registers\[4\]\[7\] rf.registers\[5\]\[7\] rf.registers\[6\]\[7\] rf.registers\[7\]\[7\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2282_ sky130_fd_sc_hd__mux4_1
X_9294_ clknet_leaf_43_clk _0454_ VGND VGND VPWR VPWR rf.registers\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8245_ _4098_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5457_ _1169_ _2194_ _2212_ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_100_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7471__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4408_ _1162_ _1163_ _1035_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8176_ net261 _3454_ _4061_ VGND VGND VPWR VPWR _4062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5700__B1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5388_ net1163 VGND VGND VPWR VPWR _2144_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7127_ net620 _3502_ _3498_ VGND VGND VPWR VPWR _3503_ sky130_fd_sc_hd__mux2_1
X_4339_ rf.registers\[28\]\[3\] rf.registers\[29\]\[3\] rf.registers\[30\]\[3\] rf.registers\[31\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__mux4_1
XANTENNA__6087__S _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7058_ _3455_ VGND VGND VPWR VPWR _3456_ sky130_fd_sc_hd__buf_4
X_6009_ _2668_ net125 _2748_ VGND VGND VPWR VPWR _2749_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_66_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4665__S1 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6550__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5090__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8477__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_57_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4656__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6460__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4690_ _1239_ _1437_ _1445_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5076__S _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4733__A1 _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6360_ net23 VGND VGND VPWR VPWR _3060_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5311_ _2065_ _2066_ _1645_ VGND VGND VPWR VPWR _2067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6291_ _3012_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8030_ _3983_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__clkbuf_1
X_5242_ _1839_ _1997_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5173_ _1927_ _1928_ _1745_ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__mux2_1
Xinput1 A1[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4344__S0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8932_ clknet_leaf_52_clk _0092_ VGND VGND VPWR VPWR rf.registers\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4944__A _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4895__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8863_ clknet_leaf_73_clk _0023_ VGND VGND VPWR VPWR rf.registers\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_7814_ _3869_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__clkbuf_1
X_8794_ clknet_leaf_17_clk _0978_ VGND VGND VPWR VPWR rf.registers\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4647__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7745_ _3069_ net1058 _3830_ VGND VGND VPWR VPWR _3833_ sky130_fd_sc_hd__mux2_1
X_4957_ _1712_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_49_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5775__A _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7466__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4888_ rf.registers\[16\]\[0\] rf.registers\[17\]\[0\] rf.registers\[18\]\[0\] rf.registers\[19\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7676_ _3796_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9415_ clknet_leaf_5_clk _0575_ VGND VGND VPWR VPWR rf.registers\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6627_ _3223_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9346_ clknet_leaf_56_clk _0506_ VGND VGND VPWR VPWR rf.registers\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6558_ net487 _3002_ _3179_ VGND VGND VPWR VPWR _3186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5509_ _2263_ _2264_ _1712_ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__mux2_1
X_9277_ clknet_leaf_15_clk _0437_ VGND VGND VPWR VPWR rf.registers\[23\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6489_ net491 _3009_ _3135_ VGND VGND VPWR VPWR _3148_ sky130_fd_sc_hd__mux2_1
X_8228_ net144 _3508_ _4083_ VGND VGND VPWR VPWR _4089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4583__S0 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8159_ _4052_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4335__S0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8154__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8000__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4574__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7417__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_85_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5860_ _2504_ _2604_ _2606_ VGND VGND VPWR VPWR _2607_ sky130_fd_sc_hd__or3_1
X_4811_ _1071_ _1566_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__nand2_1
X_5791_ _2323_ _2515_ VGND VGND VPWR VPWR _2541_ sky130_fd_sc_hd__nand2_1
XANTENNA__7286__S _3554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5595__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7530_ _3058_ net524 _3711_ VGND VGND VPWR VPWR _3719_ sky130_fd_sc_hd__mux2_1
X_4742_ _1496_ _1497_ _1259_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__mux2_1
XANTENNA__8145__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7461_ _3682_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4673_ _1254_ _1428_ _1170_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6412_ _3096_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__clkbuf_1
X_9200_ clknet_leaf_3_clk _0360_ VGND VGND VPWR VPWR rf.registers\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7392_ _3056_ net548 _3639_ VGND VGND VPWR VPWR _3646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9131_ clknet_leaf_2_clk _0291_ VGND VGND VPWR VPWR rf.registers\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6343_ _3048_ net875 _3044_ VGND VGND VPWR VPWR _3049_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9062_ clknet_leaf_0_clk _0222_ VGND VGND VPWR VPWR rf.registers\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6274_ _2254_ _2925_ _2998_ _2337_ VGND VGND VPWR VPWR _2999_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5225_ rf.registers\[20\]\[26\] rf.registers\[21\]\[26\] rf.registers\[22\]\[26\]
+ rf.registers\[23\]\[26\] _1881_ _1883_ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__mux4_1
X_8013_ _3134_ net992 _3974_ VGND VGND VPWR VPWR _3975_ sky130_fd_sc_hd__mux2_1
XANTENNA__4565__S0 _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5156_ _1908_ _1911_ _1700_ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5087_ rf.registers\[20\]\[17\] rf.registers\[21\]\[17\] rf.registers\[22\]\[17\]
+ rf.registers\[23\]\[17\] _1689_ _1693_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__mux4_1
XANTENNA__7050__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8915_ clknet_leaf_32_clk _0075_ VGND VGND VPWR VPWR rf.registers\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8846_ clknet_leaf_44_clk _0006_ VGND VGND VPWR VPWR rf.registers\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6395__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8777_ clknet_leaf_62_clk _0961_ VGND VGND VPWR VPWR rf.registers\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7196__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5989_ _2716_ _2722_ _2729_ _2621_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__o22a_1
X_7728_ _3052_ net957 _3819_ VGND VGND VPWR VPWR _3824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7659_ _3787_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7895__A0 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7924__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9329_ clknet_leaf_39_clk _0489_ VGND VGND VPWR VPWR rf.registers\[21\]\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5444__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4556__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6870__A1 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4859__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8490__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5036__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold309 rf.registers\[3\]\[18\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4795__S0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7135__A net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4547__S0 _1262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5010_ _1700_ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__buf_4
XANTENNA__6861__A1 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1009 rf.registers\[27\]\[22\] VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6074__C1 _1820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6961_ net480 _3139_ _3398_ VGND VGND VPWR VPWR _3401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8700_ clknet_leaf_16_clk _0884_ VGND VGND VPWR VPWR rf.registers\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_5912_ _2504_ _2647_ _2653_ _2656_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6892_ _3364_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8631_ clknet_leaf_33_clk _0815_ VGND VGND VPWR VPWR rf.registers\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_5843_ net81 _2102_ VGND VGND VPWR VPWR _2591_ sky130_fd_sc_hd__nor2_4
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8562_ net533 net29 _4255_ VGND VGND VPWR VPWR _4265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8118__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5774_ _2369_ _2360_ VGND VGND VPWR VPWR _2525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7513_ _3041_ net1060 _3700_ VGND VGND VPWR VPWR _3710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4725_ rf.registers\[24\]\[14\] rf.registers\[25\]\[14\] rf.registers\[26\]\[14\]
+ rf.registers\[27\]\[14\] _1324_ _1325_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_79_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8493_ _4229_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5027__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7877__A0 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4656_ rf.registers\[0\]\[7\] rf.registers\[1\]\[7\] rf.registers\[2\]\[7\] rf.registers\[3\]\[7\]
+ net120 _1193_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__mux4_1
X_7444_ _3673_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__clkbuf_1
Xhold810 rf.registers\[7\]\[19\] VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd3_1
X_7375_ _3039_ net377 _3628_ VGND VGND VPWR VPWR _3637_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold821 rf.registers\[10\]\[19\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd3_1
X_4587_ _1211_ _1342_ _1078_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__a21o_1
XANTENNA__4669__A _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5264__S _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold832 rf.registers\[26\]\[10\] VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 rf.registers\[2\]\[3\] VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9114_ clknet_leaf_37_clk _0274_ VGND VGND VPWR VPWR rf.registers\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6326_ net43 VGND VGND VPWR VPWR _3037_ sky130_fd_sc_hd__clkbuf_2
Xhold854 rf.registers\[6\]\[24\] VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 rf.registers\[16\]\[12\] VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 rf.registers\[17\]\[10\] VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 rf.registers\[28\]\[6\] VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 rf.registers\[30\]\[24\] VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4538__S0 net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6257_ net91 _2982_ VGND VGND VPWR VPWR _2983_ sky130_fd_sc_hd__xnor2_1
X_9045_ clknet_leaf_30_clk _0205_ VGND VGND VPWR VPWR rf.registers\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5208_ rf.registers\[16\]\[27\] rf.registers\[17\]\[27\] rf.registers\[18\]\[27\]
+ rf.registers\[19\]\[27\] _1767_ _1768_ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__mux4_1
X_6188_ _1978_ _2915_ VGND VGND VPWR VPWR _2917_ sky130_fd_sc_hd__nand2_1
XANTENNA__4608__S _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5139_ _1689_ VGND VGND VPWR VPWR _1895_ sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_66_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7919__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6823__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4710__S0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6368__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8829_ clknet_leaf_15_clk _1013_ VGND VGND VPWR VPWR rf.registers\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5266__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7654__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7868__A0 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5018__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4777__S0 _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8485__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5203__A _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7829__S _3843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6733__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4510_ _1260_ _1265_ _1187_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__mux2_2
X_5490_ _1671_ _2237_ _2245_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8520__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold106 rf.registers\[2\]\[26\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _1190_ _1196_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__and2_1
XANTENNA__4768__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold117 rf.registers\[5\]\[14\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold128 rf.registers\[2\]\[13\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 rf.registers\[10\]\[11\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7160_ net260 _3464_ _3517_ VGND VGND VPWR VPWR _3522_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _1087_ _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6111_ _2840_ _2844_ VGND VGND VPWR VPWR _2845_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7091_ _3478_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6042_ _2420_ _2738_ _2333_ VGND VGND VPWR VPWR _2780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5193__S0 _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5113__A _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7993_ _3964_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__clkbuf_1
X_6944_ net754 _3122_ _3387_ VGND VGND VPWR VPWR _3392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4952__A _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6875_ _3355_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7011__A1 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5248__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8614_ clknet_leaf_72_clk _0798_ VGND VGND VPWR VPWR rf.registers\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5826_ _2105_ _2573_ _2574_ _2373_ VGND VGND VPWR VPWR _2575_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5022__B1 _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6770__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5573__A1 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8545_ _4256_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__clkbuf_1
X_5757_ _2305_ _2508_ VGND VGND VPWR VPWR _2509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4708_ _1455_ _1215_ _1463_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_115_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8476_ _4220_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__clkbuf_1
X_5688_ _1926_ _2178_ VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__or2b_1
X_7427_ _3019_ net357 _3664_ VGND VGND VPWR VPWR _3665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4639_ rf.registers\[4\]\[6\] rf.registers\[5\]\[6\] rf.registers\[6\]\[6\] rf.registers\[7\]\[6\]
+ net106 _1073_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 rf.registers\[23\]\[9\] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7358_ _3627_ VGND VGND VPWR VPWR _3628_ sky130_fd_sc_hd__clkbuf_8
Xhold651 rf.registers\[31\]\[13\] VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 rf.registers\[26\]\[31\] VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 rf.registers\[10\]\[21\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlygate4sd3_1
X_6309_ _3025_ net938 _3023_ VGND VGND VPWR VPWR _3026_ sky130_fd_sc_hd__mux2_1
Xhold684 rf.registers\[6\]\[19\] VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 rf.registers\[29\]\[17\] VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6818__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7289_ _3590_ VGND VGND VPWR VPWR _3591_ sky130_fd_sc_hd__buf_4
XANTENNA__5722__S _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9028_ clknet_leaf_62_clk _0188_ VGND VGND VPWR VPWR rf.registers\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4846__B _1601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7649__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5487__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7002__A1 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7384__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8502__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5411__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6728__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5175__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output59_A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7559__S _3699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5478__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6463__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4990_ rf.registers\[12\]\[22\] rf.registers\[13\]\[22\] rf.registers\[14\]\[22\]
+ rf.registers\[15\]\[22\] _1720_ _1723_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6660_ net697 _3111_ _3231_ VGND VGND VPWR VPWR _3241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5611_ _2365_ VGND VGND VPWR VPWR _2366_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6752__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6591_ _3204_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7294__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4711__S _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8330_ net768 _3474_ _4133_ VGND VGND VPWR VPWR _4143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5542_ rf.registers\[8\]\[4\] rf.registers\[9\]\[4\] rf.registers\[10\]\[4\] rf.registers\[11\]\[4\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2298_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8261_ _4106_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5473_ _1671_ _2220_ _2224_ _2228_ VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7212_ net306 _3448_ _3539_ VGND VGND VPWR VPWR _3549_ sky130_fd_sc_hd__mux2_1
X_4424_ rf.registers\[28\]\[29\] rf.registers\[29\]\[29\] rf.registers\[30\]\[29\]
+ rf.registers\[31\]\[29\] _1173_ _1175_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8192_ net698 _3472_ _4061_ VGND VGND VPWR VPWR _4070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4355_ _1110_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__buf_4
XANTENNA__6638__S _3194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7143_ _3512_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4947__A _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7074_ net293 _3466_ _3456_ VGND VGND VPWR VPWR _3467_ sky130_fd_sc_hd__mux2_1
X_4286_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__buf_12
X_6025_ _1874_ _2743_ VGND VGND VPWR VPWR _2764_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7469__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5469__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7976_ _3955_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ net694 _3105_ _3376_ VGND VGND VPWR VPWR _3383_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6858_ _3346_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5809_ _1415_ _2557_ VGND VGND VPWR VPWR _2558_ sky130_fd_sc_hd__xor2_1
XANTENNA__6743__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9577_ clknet_leaf_6_clk _0737_ VGND VGND VPWR VPWR rf.registers\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6789_ net289 _3103_ _3304_ VGND VGND VPWR VPWR _3310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8528_ _4247_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5944__C _2160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8459_ _4211_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7932__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold470 rf.registers\[29\]\[5\] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6548__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold481 rf.registers\[8\]\[31\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5452__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold492 rf.registers\[22\]\[26\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5157__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4380__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4993__C1 _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload15 clknet_leaf_74_clk VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__clkinv_4
Xclkload26 clknet_leaf_54_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__inv_12
XFILLER_0_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload37 clknet_leaf_49_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__clkinv_4
Xclkload48 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__inv_6
Xclkload59 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload59/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5396__S0 _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5598__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4706__S _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7830_ _3877_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5320__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5776__A1 _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7761_ _3085_ net1083 _3807_ VGND VGND VPWR VPWR _3841_ sky130_fd_sc_hd__mux2_1
X_4973_ _1728_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9500_ clknet_leaf_16_clk _0660_ VGND VGND VPWR VPWR rf.registers\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6921__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6712_ _3025_ net841 _3267_ VGND VGND VPWR VPWR _3269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7692_ _3804_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9431_ clknet_leaf_23_clk _0591_ VGND VGND VPWR VPWR rf.registers\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6643_ _3232_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload9 clknet_leaf_68_clk VGND VGND VPWR VPWR clkload9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9362_ clknet_leaf_39_clk _0522_ VGND VGND VPWR VPWR rf.registers\[20\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6574_ _3019_ net928 _3195_ VGND VGND VPWR VPWR _3196_ sky130_fd_sc_hd__mux2_1
X_8313_ _4134_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5525_ _1699_ _2280_ VGND VGND VPWR VPWR _2281_ sky130_fd_sc_hd__nand2_1
X_9293_ clknet_leaf_40_clk _0453_ VGND VGND VPWR VPWR rf.registers\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8244_ _3089_ net352 _4097_ VGND VGND VPWR VPWR _4098_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5456_ _1168_ _2211_ VGND VGND VPWR VPWR _2212_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4407_ rf.registers\[0\]\[0\] rf.registers\[1\]\[0\] rf.registers\[2\]\[0\] rf.registers\[3\]\[0\]
+ net94 _1061_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__mux4_1
XANTENNA__6368__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8175_ _4060_ VGND VGND VPWR VPWR _4061_ sky130_fd_sc_hd__buf_4
XANTENNA__8149__A _4024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5387_ _1169_ _2124_ _2142_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7053__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7126_ net28 VGND VGND VPWR VPWR _3502_ sky130_fd_sc_hd__buf_2
X_4338_ _1088_ _1093_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__nand2_1
X_4269_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__buf_6
X_7057_ _3153_ _3411_ VGND VGND VPWR VPWR _3455_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_105_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6008_ _2123_ net113 _2746_ _2747_ VGND VGND VPWR VPWR _2748_ sky130_fd_sc_hd__o211a_1
XANTENNA__5301__A _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7959_ net248 _3444_ _3938_ VGND VGND VPWR VPWR _3946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6831__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6132__A _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7662__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4526__S _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5302__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7837__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6741__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8522__A _3006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7380__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5310_ rf.registers\[16\]\[2\] rf.registers\[17\]\[2\] rf.registers\[18\]\[2\] rf.registers\[19\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2066_ sky130_fd_sc_hd__mux4_1
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6290_ net824 _3011_ _3007_ VGND VGND VPWR VPWR _3012_ sky130_fd_sc_hd__mux2_1
XANTENNA__5369__S0 _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7683__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5241_ _1842_ _1996_ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_3_0__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5092__S _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5172_ rf.registers\[16\]\[29\] rf.registers\[17\]\[29\] rf.registers\[18\]\[29\]
+ rf.registers\[19\]\[29\] _1705_ _1708_ VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__mux4_1
X_8931_ clknet_leaf_52_clk _0091_ VGND VGND VPWR VPWR rf.registers\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xinput2 A1[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4344__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5541__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8862_ clknet_leaf_73_clk _0022_ VGND VGND VPWR VPWR rf.registers\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5121__A _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7813_ net342 _3502_ _3866_ VGND VGND VPWR VPWR _3869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8793_ clknet_leaf_19_clk _0977_ VGND VGND VPWR VPWR rf.registers\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7747__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4960__A _1655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7744_ _3832_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__clkbuf_1
X_4956_ _1711_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7675_ net799 _3500_ _3794_ VGND VGND VPWR VPWR _3796_ sky130_fd_sc_hd__mux2_1
XANTENNA__5267__S _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4887_ rf.registers\[20\]\[0\] rf.registers\[21\]\[0\] rf.registers\[22\]\[0\] rf.registers\[23\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9414_ clknet_leaf_5_clk _0574_ VGND VGND VPWR VPWR rf.registers\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6626_ _3075_ net447 _3217_ VGND VGND VPWR VPWR _3223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9345_ clknet_leaf_56_clk _0505_ VGND VGND VPWR VPWR rf.registers\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6557_ _3185_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5791__A _2323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5508_ rf.registers\[12\]\[6\] rf.registers\[13\]\[6\] rf.registers\[14\]\[6\] rf.registers\[15\]\[6\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_95_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9276_ clknet_leaf_16_clk _0436_ VGND VGND VPWR VPWR rf.registers\[23\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6488_ _3147_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__clkbuf_1
X_8227_ _4088_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__clkbuf_1
X_5439_ rf.registers\[24\]\[10\] rf.registers\[25\]\[10\] rf.registers\[26\]\[10\]
+ rf.registers\[27\]\[10\] _1674_ _1691_ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8158_ net1049 _3506_ _4047_ VGND VGND VPWR VPWR _4052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4583__S1 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7109_ _3490_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_8089_ _4015_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5437__B1 _2188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4335__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5177__S _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7392__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4574__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5523__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7567__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4810_ _1564_ _1565_ _1048_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__mux2_1
X_5790_ _2271_ _2538_ VGND VGND VPWR VPWR _2540_ sky130_fd_sc_hd__nor2_1
X_4741_ rf.registers\[16\]\[15\] rf.registers\[17\]\[15\] rf.registers\[18\]\[15\]
+ rf.registers\[19\]\[15\] net128 _1263_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7460_ _3056_ net1132 _3675_ VGND VGND VPWR VPWR _3682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4672_ _1426_ _1427_ _1211_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__mux2_1
X_6411_ net800 _3095_ _3093_ VGND VGND VPWR VPWR _3096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8398__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7391_ _3645_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9130_ clknet_leaf_45_clk _0290_ VGND VGND VPWR VPWR rf.registers\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6342_ net17 VGND VGND VPWR VPWR _3048_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9061_ clknet_leaf_57_clk _0221_ VGND VGND VPWR VPWR rf.registers\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6273_ _2958_ _2997_ _2363_ VGND VGND VPWR VPWR _2998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8012_ _3951_ VGND VGND VPWR VPWR _3974_ sky130_fd_sc_hd__clkbuf_8
X_5224_ _1800_ _1979_ VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4955__A net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6646__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5155_ _1909_ _1910_ _1745_ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__mux2_1
XANTENNA__7331__A _3590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5086_ _1638_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_108_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8914_ clknet_leaf_25_clk _0074_ VGND VGND VPWR VPWR rf.registers\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4642__B2 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8845_ clknet_leaf_43_clk _0005_ VGND VGND VPWR VPWR rf.registers\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7477__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5786__A _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8776_ clknet_leaf_63_clk _0960_ VGND VGND VPWR VPWR rf.registers\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7592__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5988_ net123 _2728_ VGND VGND VPWR VPWR _2729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7727_ _3823_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__clkbuf_1
X_4939_ _1688_ _1694_ _1686_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7658_ net210 _3483_ _3783_ VGND VGND VPWR VPWR _3787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6609_ _3058_ net340 _3206_ VGND VGND VPWR VPWR _3214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7589_ _3750_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
X_9328_ clknet_leaf_13_clk _0488_ VGND VGND VPWR VPWR rf.registers\[21\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6410__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9259_ clknet_leaf_2_clk _0419_ VGND VGND VPWR VPWR rf.registers\[23\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7940__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5658__B1 _2097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5026__A _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4556__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6556__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5460__S _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5696__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5635__S _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6320__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4795__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4547__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6466__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7151__A _3516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8063__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6960_ _3400_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_37_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5911_ _2654_ _2655_ VGND VGND VPWR VPWR _2656_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6891_ net595 _3137_ _3362_ VGND VGND VPWR VPWR _3364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4714__S _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8630_ clknet_leaf_24_clk _0814_ VGND VGND VPWR VPWR rf.registers\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_5842_ _1666_ _2040_ VGND VGND VPWR VPWR _2590_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8561_ _4264_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5773_ _2338_ _2365_ VGND VGND VPWR VPWR _2524_ sky130_fd_sc_hd__nor2_1
XANTENNA__6214__B _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7512_ _3709_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
X_4724_ _1215_ _1471_ _1475_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__a2bb2o_2
X_8492_ net536 net27 _4227_ VGND VGND VPWR VPWR _4229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7443_ _3039_ net747 _3664_ VGND VGND VPWR VPWR _3673_ sky130_fd_sc_hd__mux2_1
X_4655_ rf.registers\[4\]\[7\] rf.registers\[5\]\[7\] rf.registers\[6\]\[7\] rf.registers\[7\]\[7\]
+ net120 _1193_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold800 rf.registers\[26\]\[22\] VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd3_1
X_7374_ _3636_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold811 rf.registers\[18\]\[29\] VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4586_ rf.registers\[8\]\[30\] rf.registers\[9\]\[30\] rf.registers\[10\]\[30\] rf.registers\[11\]\[30\]
+ net135 _1184_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__mux4_1
Xhold822 rf.registers\[11\]\[28\] VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 rf.registers\[23\]\[31\] VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlygate4sd3_1
X_9113_ clknet_leaf_19_clk _0273_ VGND VGND VPWR VPWR rf.registers\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold844 rf.registers\[31\]\[25\] VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd3_1
X_6325_ _3036_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__clkbuf_1
Xhold855 rf.registers\[4\]\[24\] VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold866 rf.registers\[1\]\[21\] VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold877 rf.registers\[0\]\[28\] VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 rf.registers\[15\]\[1\] VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__dlygate4sd3_1
X_9044_ clknet_leaf_30_clk _0204_ VGND VGND VPWR VPWR rf.registers\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold899 rf.registers\[27\]\[11\] VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ _2741_ _2981_ VGND VGND VPWR VPWR _2982_ sky130_fd_sc_hd__nor2_1
XANTENNA__4538__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5207_ rf.registers\[20\]\[27\] rf.registers\[21\]\[27\] rf.registers\[22\]\[27\]
+ rf.registers\[23\]\[27\] _1767_ _1768_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__mux4_1
X_6187_ _1978_ _2915_ VGND VGND VPWR VPWR _2916_ sky130_fd_sc_hd__or2_1
XANTENNA__7061__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8054__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5138_ _1773_ _1893_ VGND VGND VPWR VPWR _1894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5069_ rf.registers\[28\]\[19\] rf.registers\[29\]\[19\] rf.registers\[30\]\[19\]
+ rf.registers\[31\]\[19\] _1676_ _1681_ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__mux4_1
XANTENNA__4710__S1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8828_ clknet_leaf_16_clk _1012_ VGND VGND VPWR VPWR rf.registers\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7000__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8759_ clknet_leaf_24_clk _0943_ VGND VGND VPWR VPWR rf.registers\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4777__S1 _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7670__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4595__A _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5203__B _1958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8006__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7845__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5365__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4440_ rf.registers\[12\]\[29\] rf.registers\[13\]\[29\] rf.registers\[14\]\[29\]
+ rf.registers\[15\]\[29\] _1192_ _1195_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__mux4_1
XANTENNA__6531__A1 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold107 rf.registers\[1\]\[17\] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4768__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold118 rf.registers\[5\]\[10\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 rf.registers\[5\]\[1\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4371_ _1111_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__and2_2
X_6110_ _2827_ _2831_ _2843_ VGND VGND VPWR VPWR _2844_ sky130_fd_sc_hd__a21boi_1
X_7090_ net1081 _3476_ _3477_ VGND VGND VPWR VPWR _3478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6041_ _2704_ _2778_ _1879_ VGND VGND VPWR VPWR _2779_ sky130_fd_sc_hd__mux2_1
XANTENNA__6196__S _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5193__S1 _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7992_ _3113_ net778 _3963_ VGND VGND VPWR VPWR _3964_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9152__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6943_ _3391_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7547__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6874_ net202 _3120_ _3351_ VGND VGND VPWR VPWR _3355_ sky130_fd_sc_hd__mux2_1
XANTENNA__6225__A _1942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8613_ clknet_leaf_52_clk _0797_ VGND VGND VPWR VPWR rf.registers\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5825_ _2255_ _2461_ _2463_ _2337_ VGND VGND VPWR VPWR _2574_ sky130_fd_sc_hd__o22a_1
XANTENNA__5022__A1 _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7755__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8544_ net308 net19 _4255_ VGND VGND VPWR VPWR _4256_ sky130_fd_sc_hd__mux2_1
X_5756_ _1060_ _2507_ VGND VGND VPWR VPWR _2508_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4781__B1 _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4707_ _1457_ _1459_ _1462_ _1071_ _1057_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8475_ net230 net18 _4216_ VGND VGND VPWR VPWR _4220_ sky130_fd_sc_hd__mux2_1
XANTENNA__5275__S _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5687_ _2252_ _2437_ _2440_ VGND VGND VPWR VPWR _2441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7056__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7426_ _3663_ VGND VGND VPWR VPWR _3664_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6522__A1 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4638_ _1036_ _1393_ _1037_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold630 rf.registers\[16\]\[23\] VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd3_1
X_7357_ _3020_ _3626_ VGND VGND VPWR VPWR _3627_ sky130_fd_sc_hd__nand2_4
Xhold641 rf.registers\[20\]\[6\] VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _1029_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold652 rf.registers\[21\]\[22\] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold663 rf.registers\[0\]\[27\] VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ net25 VGND VGND VPWR VPWR _3025_ sky130_fd_sc_hd__clkbuf_2
Xhold674 rf.registers\[30\]\[26\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 rf.registers\[23\]\[23\] VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7288_ _3193_ _3553_ VGND VGND VPWR VPWR _3590_ sky130_fd_sc_hd__nand2_4
Xhold696 rf.registers\[21\]\[10\] VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd3_1
X_9027_ clknet_leaf_67_clk _0187_ VGND VGND VPWR VPWR rf.registers\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6239_ _2965_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8496__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4529__S _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5907__A1_N _2458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5175__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6029__B1 _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4686__S0 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4460__C1 _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7575__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5610_ _1169_ _2098_ _1803_ VGND VGND VPWR VPWR _2365_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6590_ _3039_ net532 _3195_ VGND VGND VPWR VPWR _3204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5541_ rf.registers\[12\]\[4\] rf.registers\[13\]\[4\] rf.registers\[14\]\[4\] rf.registers\[15\]\[4\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_65_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8260_ _3109_ net279 _4097_ VGND VGND VPWR VPWR _4106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5472_ _1717_ _2227_ _1729_ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__a21oi_1
X_7211_ _3548_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4423_ _1176_ _1177_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__mux2_1
XANTENNA__6919__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8191_ _4069_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7604__A _3735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7142_ net396 _3446_ _3498_ VGND VGND VPWR VPWR _3512_ sky130_fd_sc_hd__mux2_1
X_4354_ _1057_ _1094_ _1098_ _1102_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a32o_2
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7073_ net41 VGND VGND VPWR VPWR _3466_ sky130_fd_sc_hd__buf_2
X_4285_ A2[0] VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__buf_12
X_6024_ _1858_ _2762_ VGND VGND VPWR VPWR _2763_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6654__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4963__A _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7975_ _3097_ net985 _3952_ VGND VGND VPWR VPWR _3955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6926_ _3382_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6857_ net334 _3103_ _3340_ VGND VGND VPWR VPWR _3346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7485__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4429__S0 _1182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4902__S _1645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5808_ net118 net95 net131 _2411_ VGND VGND VPWR VPWR _2557_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9576_ clknet_leaf_65_clk _0736_ VGND VGND VPWR VPWR rf.registers\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6788_ _3309_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8527_ net701 net42 _4244_ VGND VGND VPWR VPWR _4247_ sky130_fd_sc_hd__mux2_1
XANTENNA__4754__B1 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5739_ _2490_ _2179_ _2426_ VGND VGND VPWR VPWR _2491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8458_ net267 net41 _4205_ VGND VGND VPWR VPWR _4211_ sky130_fd_sc_hd__mux2_1
XANTENNA__8496__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7409_ _3073_ net876 _3650_ VGND VGND VPWR VPWR _3655_ sky130_fd_sc_hd__mux2_1
XANTENNA__6829__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8389_ _4174_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4601__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold460 rf.registers\[24\]\[4\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 rf.registers\[15\]\[12\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 rf.registers\[14\]\[0\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 rf.registers\[14\]\[18\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5157__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6564__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7759__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4873__A _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload16 clknet_leaf_1_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload27 clknet_leaf_55_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8487__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload38 clknet_leaf_50_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_134_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload49 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload49/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6739__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5396__S1 _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output71_A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7998__A0 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8411__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7760_ _3840_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__clkbuf_1
X_4972_ net5 VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__buf_4
XANTENNA__6973__A1 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5320__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6711_ _3268_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_82_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7691_ net571 _3448_ _3794_ VGND VGND VPWR VPWR _3804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9430_ clknet_leaf_24_clk _0590_ VGND VGND VPWR VPWR rf.registers\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6642_ net219 _3089_ _3231_ VGND VGND VPWR VPWR _3232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4722__S _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6503__A _3156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9361_ clknet_leaf_39_clk _0521_ VGND VGND VPWR VPWR rf.registers\[20\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6573_ _3194_ VGND VGND VPWR VPWR _3195_ sky130_fd_sc_hd__buf_4
XFILLER_0_143_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8312_ net258 _3454_ _4133_ VGND VGND VPWR VPWR _4134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5524_ _2278_ _2279_ _1685_ VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9292_ clknet_leaf_50_clk _0452_ VGND VGND VPWR VPWR rf.registers\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8243_ _4096_ VGND VGND VPWR VPWR _4097_ sky130_fd_sc_hd__buf_4
X_5455_ _1639_ _2210_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4406_ rf.registers\[4\]\[0\] rf.registers\[5\]\[0\] rf.registers\[6\]\[0\] rf.registers\[7\]\[0\]
+ net94 _1061_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8174_ _3091_ _3153_ VGND VGND VPWR VPWR _4060_ sky130_fd_sc_hd__nor2_4
X_5386_ _1669_ _2141_ VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7125_ _3501_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
X_4337_ _1091_ _1092_ _1040_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__mux2_1
XANTENNA__7989__A0 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7056_ net14 VGND VGND VPWR VPWR _3454_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4268_ net8 VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6007_ _2123_ net113 _2726_ VGND VGND VPWR VPWR _2747_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7958_ _3945_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6909_ net790 _3015_ _3339_ VGND VGND VPWR VPWR _3373_ sky130_fd_sc_hd__mux2_1
X_7889_ _3002_ net731 _3902_ VGND VGND VPWR VPWR _3909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6413__A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8104__S _3988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5075__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6132__B _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9559_ clknet_leaf_26_clk _0719_ VGND VGND VPWR VPWR rf.registers\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4822__S0 _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8469__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5463__S _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold290 rf.registers\[27\]\[13\] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5302__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6323__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7853__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4813__S0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5881__B _2626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5369__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5240_ _1777_ _1987_ _1995_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__a21oi_4
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5171_ rf.registers\[20\]\[29\] rf.registers\[21\]\[29\] rf.registers\[22\]\[29\]
+ rf.registers\[23\]\[29\] _1705_ _1708_ VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8930_ clknet_leaf_56_clk _0090_ VGND VGND VPWR VPWR rf.registers\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xinput3 A1[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5541__S1 _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8861_ clknet_leaf_16_clk _0021_ VGND VGND VPWR VPWR rf.registers\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_7812_ _3868_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__clkbuf_1
X_8792_ clknet_leaf_27_clk _0976_ VGND VGND VPWR VPWR rf.registers\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7743_ _3067_ net1067 _3830_ VGND VGND VPWR VPWR _3832_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4955_ net3 VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7674_ _3795_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_1
X_4886_ net2 VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5057__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9413_ clknet_leaf_54_clk _0573_ VGND VGND VPWR VPWR rf.registers\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6625_ _3222_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7763__S _3807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4804__S0 _1042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6556_ net588 _3145_ _3179_ VGND VGND VPWR VPWR _3185_ sky130_fd_sc_hd__mux2_1
X_9344_ clknet_leaf_60_clk _0504_ VGND VGND VPWR VPWR rf.registers\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5507_ rf.registers\[8\]\[6\] rf.registers\[9\]\[6\] rf.registers\[10\]\[6\] rf.registers\[11\]\[6\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2263_ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9275_ clknet_leaf_34_clk _0435_ VGND VGND VPWR VPWR rf.registers\[23\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6487_ net688 _3002_ _3135_ VGND VGND VPWR VPWR _3147_ sky130_fd_sc_hd__mux2_1
XANTENNA__7064__A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8226_ net497 _3506_ _4083_ VGND VGND VPWR VPWR _4088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5438_ _2144_ _2193_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5685__A1 _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8157_ _4051_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__clkbuf_1
X_5369_ rf.registers\[20\]\[14\] rf.registers\[21\]\[14\] rf.registers\[22\]\[14\]
+ rf.registers\[23\]\[14\] _1733_ _1679_ VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__mux4_1
X_7108_ net427 _3489_ _3477_ VGND VGND VPWR VPWR _3490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8088_ net696 _3504_ _4011_ VGND VGND VPWR VPWR _4015_ sky130_fd_sc_hd__mux2_1
XANTENNA__6634__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5437__A1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7039_ net621 _3442_ _3435_ VGND VGND VPWR VPWR _3443_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7938__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6143__A _2033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7673__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7114__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5523__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6752__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_124_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5287__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4740_ rf.registers\[20\]\[15\] rf.registers\[21\]\[15\] rf.registers\[22\]\[15\]
+ rf.registers\[23\]\[15\] net128 _1263_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5039__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4671_ rf.registers\[0\]\[23\] rf.registers\[1\]\[23\] rf.registers\[2\]\[23\] rf.registers\[3\]\[23\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6410_ net25 VGND VGND VPWR VPWR _3095_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7390_ _3054_ net1071 _3639_ VGND VGND VPWR VPWR _3645_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6341_ _3047_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8302__A0 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7105__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9060_ clknet_leaf_62_clk _0220_ VGND VGND VPWR VPWR rf.registers\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4301__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6272_ _2379_ _2377_ VGND VGND VPWR VPWR _2997_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5211__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8011_ _3973_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5223_ _1842_ _1978_ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__nor2_1
XANTENNA__6927__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5154_ rf.registers\[24\]\[30\] rf.registers\[25\]\[30\] rf.registers\[26\]\[30\]
+ rf.registers\[27\]\[30\] _1895_ _1897_ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__mux4_1
XANTENNA__6616__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5085_ _1669_ _1821_ _1840_ VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8913_ clknet_leaf_42_clk _0073_ VGND VGND VPWR VPWR rf.registers\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_142_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8844_ clknet_leaf_46_clk _0004_ VGND VGND VPWR VPWR rf.registers\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5187__A_N net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8775_ clknet_leaf_2_clk _0959_ VGND VGND VPWR VPWR rf.registers\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5987_ _2726_ _2727_ VGND VGND VPWR VPWR _2728_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_121_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7726_ _3050_ net933 _3819_ VGND VGND VPWR VPWR _3823_ sky130_fd_sc_hd__mux2_1
X_4938_ rf.registers\[24\]\[23\] rf.registers\[25\]\[23\] rf.registers\[26\]\[23\]
+ rf.registers\[27\]\[23\] _1689_ _1693_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7657_ _3786_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__clkbuf_1
X_4869_ _1621_ _1624_ _1213_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6608_ _3213_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__clkbuf_1
X_7588_ _3048_ net1013 _3747_ VGND VGND VPWR VPWR _3750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5450__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9327_ clknet_leaf_10_clk _0487_ VGND VGND VPWR VPWR rf.registers\[21\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6539_ net658 _3128_ _3168_ VGND VGND VPWR VPWR _3176_ sky130_fd_sc_hd__mux2_1
XANTENNA__5307__A _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9258_ clknet_leaf_8_clk _0418_ VGND VGND VPWR VPWR rf.registers\[23\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8209_ net488 _3489_ _4072_ VGND VGND VPWR VPWR _4079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6837__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9189_ clknet_leaf_61_clk _0349_ VGND VGND VPWR VPWR rf.registers\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6607__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6138__A _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7280__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7668__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8353__A _4132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5269__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5696__B _1660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5594__B1 _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5217__A _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6747__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5651__S _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6048__A _1820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6482__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5910_ _2471_ _2605_ _2591_ _2462_ VGND VGND VPWR VPWR _2655_ sky130_fd_sc_hd__a22o_1
X_6890_ _3363_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5841_ _1880_ _2588_ _2421_ VGND VGND VPWR VPWR _2589_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5772_ _1111_ _2522_ _2487_ _2382_ VGND VGND VPWR VPWR _2523_ sky130_fd_sc_hd__o2bb2a_1
X_8560_ net599 net28 _4255_ VGND VGND VPWR VPWR _4264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7511_ _3039_ net666 _3700_ VGND VGND VPWR VPWR _3709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4723_ _1205_ _1478_ _1170_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8491_ _4228_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7442_ _3672_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4654_ _1071_ _1409_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5888__A1 _2229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5888__B2 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7373_ _3037_ net886 _3628_ VGND VGND VPWR VPWR _3636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold801 rf.registers\[13\]\[6\] VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6230__B _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4585_ _1189_ _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__and2_1
Xhold812 rf.registers\[28\]\[3\] VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5127__A _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold823 rf.registers\[22\]\[7\] VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6324_ _3035_ net1038 _3023_ VGND VGND VPWR VPWR _3036_ sky130_fd_sc_hd__mux2_1
Xhold834 rf.registers\[22\]\[14\] VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd3_1
X_9112_ clknet_leaf_11_clk _0272_ VGND VGND VPWR VPWR rf.registers\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold845 rf.registers\[21\]\[9\] VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold856 rf.registers\[22\]\[1\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 rf.registers\[29\]\[10\] VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 rf.registers\[13\]\[20\] VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__dlygate4sd3_1
X_9043_ clknet_leaf_34_clk _0203_ VGND VGND VPWR VPWR rf.registers\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6255_ net1157 _2929_ VGND VGND VPWR VPWR _2981_ sky130_fd_sc_hd__nor2_1
Xhold889 rf.registers\[26\]\[20\] VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4966__A _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5561__S _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5206_ _1926_ _1961_ _1877_ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__mux2_1
X_6186_ net99 _2914_ VGND VGND VPWR VPWR _2915_ sky130_fd_sc_hd__xor2_1
X_5137_ _1891_ _1892_ _1889_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_150_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5068_ rf.registers\[24\]\[19\] rf.registers\[25\]\[19\] rf.registers\[26\]\[19\]
+ rf.registers\[27\]\[19\] _1822_ _1823_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__mux4_1
XANTENNA__6392__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8827_ clknet_leaf_22_clk _1011_ VGND VGND VPWR VPWR rf.registers\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8758_ clknet_leaf_25_clk _0942_ VGND VGND VPWR VPWR rf.registers\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7709_ _3033_ net1136 _3808_ VGND VGND VPWR VPWR _3814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8689_ clknet_leaf_29_clk _0873_ VGND VGND VPWR VPWR rf.registers\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8112__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7951__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5471__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4303__A1 _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7253__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7398__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4550__S _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5319__B1 _1655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold108 rf.registers\[17\]\[15\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold119 rf.registers\[6\]\[4\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ net85 VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6040_ _2734_ _2777_ _1877_ VGND VGND VPWR VPWR _2778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7991_ _3951_ VGND VGND VPWR VPWR _3963_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6942_ net225 _3120_ _3387_ VGND VGND VPWR VPWR _3391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6873_ _3354_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8612_ clknet_leaf_52_clk _0796_ VGND VGND VPWR VPWR rf.registers\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6940__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ _2470_ _2460_ _2252_ VGND VGND VPWR VPWR _2573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5755_ _2411_ net95 VGND VGND VPWR VPWR _2507_ sky130_fd_sc_hd__nor2_1
X_8543_ _3006_ VGND VGND VPWR VPWR _4255_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4781__A1 _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4706_ _1460_ _1461_ _1048_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8474_ _4219_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__clkbuf_1
X_5686_ _2252_ _2439_ VGND VGND VPWR VPWR _2440_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7425_ _3552_ _3626_ VGND VGND VPWR VPWR _3663_ sky130_fd_sc_hd__nand2_4
X_4637_ rf.registers\[12\]\[6\] rf.registers\[13\]\[6\] rf.registers\[14\]\[6\] rf.registers\[15\]\[6\]
+ net120 _1193_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7771__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold620 rf.registers\[4\]\[20\] VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__dlygate4sd3_1
X_7356_ net11 net12 net13 VGND VGND VPWR VPWR _3626_ sky130_fd_sc_hd__and3b_2
X_4568_ _1027_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__clkbuf_8
Xhold631 rf.registers\[23\]\[22\] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 rf.registers\[14\]\[28\] VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold653 rf.registers\[8\]\[16\] VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd3_1
X_6307_ _3024_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__clkbuf_1
Xhold664 rf.registers\[23\]\[18\] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__dlygate4sd3_1
X_7287_ _3589_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
Xhold675 rf.registers\[16\]\[27\] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 rf.registers\[16\]\[9\] VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd3_1
X_4499_ _1248_ _1250_ _1253_ _1254_ _1170_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__a221o_1
Xhold697 rf.registers\[30\]\[1\] VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__dlygate4sd3_1
X_9026_ clknet_leaf_59_clk _0186_ VGND VGND VPWR VPWR rf.registers\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6238_ _2964_ _2957_ _2963_ VGND VGND VPWR VPWR _2965_ sky130_fd_sc_hd__or3_4
X_6169_ _2613_ _2737_ _2898_ _2899_ VGND VGND VPWR VPWR _2900_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6416__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7011__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone20 net108 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_16
Xclone53 _1181_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_20_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7681__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6277__A1 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7777__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8017__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6326__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4686__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7856__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6760__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5540_ _2292_ _2295_ _1696_ VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6061__A _2737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5471_ _2225_ _2226_ _1739_ VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4422_ _1036_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__buf_4
X_7210_ net359 _3446_ _3539_ VGND VGND VPWR VPWR _3548_ sky130_fd_sc_hd__mux2_1
X_8190_ net983 _3470_ _4061_ VGND VGND VPWR VPWR _4069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7141_ _3511_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
X_4353_ _1108_ _1088_ net8 VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7072_ _3465_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
X_4284_ _1034_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__buf_4
X_6023_ _1601_ _2761_ VGND VGND VPWR VPWR _2762_ sky130_fd_sc_hd__xor2_1
XANTENNA__4374__S0 _1065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7974_ _3954_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5140__A _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6925_ net1088 _3103_ _3376_ VGND VGND VPWR VPWR _3382_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6856_ _3345_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4429__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5807_ _2504_ _2544_ _2545_ _2556_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__a31o_4
X_9575_ clknet_leaf_5_clk _0735_ VGND VGND VPWR VPWR rf.registers\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6787_ net201 _3101_ _3304_ VGND VGND VPWR VPWR _3309_ sky130_fd_sc_hd__mux2_1
XANTENNA__7940__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8987__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7067__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8526_ _4246_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4754__A1 _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5951__B1 _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5738_ _1878_ VGND VGND VPWR VPWR _2490_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8457_ _4210_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__clkbuf_1
X_5669_ _1876_ VGND VGND VPWR VPWR _2423_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7408_ _3654_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8388_ net619 _3464_ _4169_ VGND VGND VPWR VPWR _4174_ sky130_fd_sc_hd__mux2_1
XANTENNA__4601__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold450 rf.registers\[15\]\[8\] VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 rf.registers\[3\]\[24\] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
X_7339_ _3617_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
Xhold472 rf.registers\[2\]\[23\] VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7456__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold483 rf.registers\[12\]\[29\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 rf.registers\[12\]\[27\] VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9009_ clknet_leaf_41_clk _0169_ VGND VGND VPWR VPWR rf.registers\[31\]\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4365__S0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_51_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6580__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4993__A1 _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8184__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload17 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload17/X sky130_fd_sc_hd__clkbuf_4
Xclkload28 clknet_leaf_56_clk VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__inv_6
XFILLER_0_63_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload39 clknet_leaf_51_clk VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8300__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5170__A1 _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output64_A net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4356__S0 _1042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6056__A _2458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4971_ _1724_ _1725_ _1726_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__mux2_1
XANTENNA__7586__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6710_ _3019_ net564 _3267_ VGND VGND VPWR VPWR _3268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7690_ _3803_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6641_ _3230_ VGND VGND VPWR VPWR _3231_ sky130_fd_sc_hd__buf_4
XFILLER_0_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4304__A _1059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9360_ clknet_leaf_13_clk _0520_ VGND VGND VPWR VPWR rf.registers\[20\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6572_ _3192_ _3193_ VGND VGND VPWR VPWR _3194_ sky130_fd_sc_hd__nand2_4
XFILLER_0_144_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8311_ _4132_ VGND VGND VPWR VPWR _4133_ sky130_fd_sc_hd__clkbuf_8
X_5523_ rf.registers\[8\]\[7\] rf.registers\[9\]\[7\] rf.registers\[10\]\[7\] rf.registers\[11\]\[7\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__mux4_1
X_9291_ clknet_leaf_1_clk _0451_ VGND VGND VPWR VPWR rf.registers\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8242_ _3552_ _3192_ VGND VGND VPWR VPWR _4096_ sky130_fd_sc_hd__nand2_4
X_5454_ _1670_ _2201_ _2205_ _2209_ VGND VGND VPWR VPWR _2210_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4405_ _1038_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5385_ _1639_ _2140_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__nor2_1
X_8173_ _4059_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4336_ rf.registers\[16\]\[3\] rf.registers\[17\]\[3\] rf.registers\[18\]\[3\] rf.registers\[19\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__mux4_1
X_7124_ net706 _3500_ _3498_ VGND VGND VPWR VPWR _3501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4347__S0 _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6665__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7055_ _3453_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6006_ net110 _2713_ _2725_ VGND VGND VPWR VPWR _2746_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_19_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7957_ net650 _3442_ _3938_ VGND VGND VPWR VPWR _3945_ sky130_fd_sc_hd__mux2_1
XANTENNA__5621__C1 _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6908_ _3372_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8166__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7888_ _3908_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6839_ net592 _3013_ _3326_ VGND VGND VPWR VPWR _3336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7913__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5075__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9558_ clknet_leaf_25_clk _0718_ VGND VGND VPWR VPWR rf.registers\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4822__S1 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8509_ _4237_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9489_ clknet_leaf_39_clk _0649_ VGND VGND VPWR VPWR rf.registers\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8120__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4586__S0 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold280 rf.registers\[0\]\[4\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 rf.registers\[9\]\[3\] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4884__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6652__A1 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6168__B1 _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4813__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6340__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6891__A1 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5170_ _1169_ _1905_ _1925_ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6485__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 A1[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
X_8860_ clknet_leaf_18_clk _0020_ VGND VGND VPWR VPWR rf.registers\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7811_ net740 _3500_ _3866_ VGND VGND VPWR VPWR _3868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8791_ clknet_leaf_23_clk _0975_ VGND VGND VPWR VPWR rf.registers\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8205__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7742_ _3831_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4501__S0 _1220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4954_ rf.registers\[12\]\[23\] rf.registers\[13\]\[23\] rf.registers\[14\]\[23\]
+ rf.registers\[15\]\[23\] _1705_ _1708_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7673_ net714 _3497_ _3794_ VGND VGND VPWR VPWR _3795_ sky130_fd_sc_hd__mux2_1
X_4885_ net1 VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9412_ clknet_leaf_51_clk _0572_ VGND VGND VPWR VPWR rf.registers\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5057__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6624_ _3073_ net776 _3217_ VGND VGND VPWR VPWR _3222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4804__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9343_ clknet_leaf_73_clk _0503_ VGND VGND VPWR VPWR rf.registers\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6555_ _3184_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5506_ _2258_ _2261_ _1696_ VGND VGND VPWR VPWR _2262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9274_ clknet_leaf_35_clk _0434_ VGND VGND VPWR VPWR rf.registers\[23\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8320__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6486_ _3146_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__clkbuf_1
X_8225_ _4087_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__clkbuf_1
X_5437_ _1670_ _2184_ _2188_ _2192_ VGND VGND VPWR VPWR _2193_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5368_ _1639_ _2123_ VGND VGND VPWR VPWR _2124_ sky130_fd_sc_hd__nor2_1
X_8156_ net160 _3504_ _4047_ VGND VGND VPWR VPWR _4051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6395__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7107_ net21 VGND VGND VPWR VPWR _3489_ sky130_fd_sc_hd__buf_2
X_4319_ rf.registers\[12\]\[5\] rf.registers\[13\]\[5\] rf.registers\[14\]\[5\] rf.registers\[15\]\[5\]
+ net106 _1073_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__mux4_1
X_5299_ rf.registers\[12\]\[3\] rf.registers\[13\]\[3\] rf.registers\[14\]\[3\] rf.registers\[15\]\[3\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__mux4_1
X_8087_ _4014_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__clkbuf_1
X_7038_ net32 VGND VGND VPWR VPWR _3442_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4740__S0 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8989_ clknet_leaf_3_clk _0149_ VGND VGND VPWR VPWR rf.registers\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8139__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload9_A clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4553__S _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5287__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8025__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7864__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5039__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4670_ rf.registers\[4\]\[23\] rf.registers\[5\]\[23\] rf.registers\[6\]\[23\] rf.registers\[7\]\[23\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8550__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4798__S0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6340_ _3046_ net1075 _3044_ VGND VGND VPWR VPWR _3047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6271_ _2942_ VGND VGND VPWR VPWR _2996_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5211__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8010_ _3132_ net1116 _3963_ VGND VGND VPWR VPWR _3973_ sky130_fd_sc_hd__mux2_1
X_5222_ _1777_ _1969_ _1973_ _1977_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_90_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5153_ rf.registers\[28\]\[30\] rf.registers\[29\]\[30\] rf.registers\[30\]\[30\]
+ rf.registers\[31\]\[30\] _1895_ _1897_ VGND VGND VPWR VPWR _1909_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_90_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5084_ _1758_ _1838_ _1839_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__o21a_1
XANTENNA__4627__B1 _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8912_ clknet_leaf_12_clk _0072_ VGND VGND VPWR VPWR rf.registers\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8843_ clknet_leaf_4_clk _0003_ VGND VGND VPWR VPWR rf.registers\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8774_ clknet_leaf_2_clk _0958_ VGND VGND VPWR VPWR rf.registers\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5986_ net110 _2714_ VGND VGND VPWR VPWR _2727_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_121_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7725_ _3822_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4937_ _1692_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 _3412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7656_ net161 _3481_ _3783_ VGND VGND VPWR VPWR _3786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4868_ _1622_ _1623_ _1259_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__mux2_1
XANTENNA__8541__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6607_ _3056_ net934 _3206_ VGND VGND VPWR VPWR _3213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7587_ _3749_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
X_4799_ rf.registers\[0\]\[10\] rf.registers\[1\]\[10\] rf.registers\[2\]\[10\] rf.registers\[3\]\[10\]
+ net107 _1105_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5450__S1 _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9326_ clknet_leaf_41_clk _0486_ VGND VGND VPWR VPWR rf.registers\[21\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6538_ _3175_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5307__B _2062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9257_ clknet_leaf_49_clk _0417_ VGND VGND VPWR VPWR rf.registers\[23\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6469_ _3092_ VGND VGND VPWR VPWR _3135_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6855__A1 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8208_ _4078_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__clkbuf_1
X_9188_ clknet_leaf_62_clk _0348_ VGND VGND VPWR VPWR rf.registers\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8139_ net663 _3487_ _4036_ VGND VGND VPWR VPWR _4042_ sky130_fd_sc_hd__mux2_1
XANTENNA__6419__A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7949__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6853__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4713__S0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5269__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8296__A0 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4999__A_N _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4857__B1 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6329__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4704__S0 net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7023__A1 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5840_ _2040_ _2372_ VGND VGND VPWR VPWR _2588_ sky130_fd_sc_hd__nand2_2
XFILLER_0_76_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5771_ _2388_ _2397_ _1126_ VGND VGND VPWR VPWR _2522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7594__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7510_ _3708_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4722_ _1476_ _1477_ _1198_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8490_ net268 net26 _4227_ VGND VGND VPWR VPWR _4228_ sky130_fd_sc_hd__mux2_1
XANTENNA__8523__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7441_ _3037_ net659 _3664_ VGND VGND VPWR VPWR _3672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4653_ _1407_ _1408_ _1040_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput40 WD3[4] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XFILLER_0_114_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7372_ _3635_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
X_4584_ rf.registers\[12\]\[30\] rf.registers\[13\]\[30\] rf.registers\[14\]\[30\]
+ rf.registers\[15\]\[30\] net127 _1222_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__mux4_1
Xhold802 rf.registers\[15\]\[22\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold813 rf.registers\[12\]\[16\] VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd3_1
X_9111_ clknet_leaf_33_clk _0271_ VGND VGND VPWR VPWR rf.registers\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6323_ net42 VGND VGND VPWR VPWR _3035_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_92_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold824 rf.registers\[17\]\[30\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6938__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold835 rf.registers\[10\]\[20\] VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 rf.registers\[15\]\[0\] VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 rf.registers\[8\]\[19\] VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6837__A1 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold868 rf.registers\[22\]\[15\] VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__dlygate4sd3_1
X_9042_ clknet_leaf_39_clk _0202_ VGND VGND VPWR VPWR rf.registers\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5196__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6254_ _2974_ _2797_ _2979_ _2421_ VGND VGND VPWR VPWR _2980_ sky130_fd_sc_hd__o211a_1
Xhold879 rf.registers\[31\]\[30\] VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5205_ _1944_ _1960_ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__or2_1
X_6185_ _1447_ _1299_ _2901_ _2871_ _2741_ VGND VGND VPWR VPWR _2914_ sky130_fd_sc_hd__a41o_1
XANTENNA__6239__A _2965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5136_ rf.registers\[12\]\[31\] rf.registers\[13\]\[31\] rf.registers\[14\]\[31\]
+ rf.registers\[15\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7769__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4982__A _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6673__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5067_ _1735_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_123_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5289__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8826_ clknet_leaf_20_clk _1010_ VGND VGND VPWR VPWR rf.registers\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6405__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8757_ clknet_leaf_32_clk _0941_ VGND VGND VPWR VPWR rf.registers\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_5969_ _2710_ _1494_ VGND VGND VPWR VPWR _2711_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_43_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7708_ _3813_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_101_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8688_ clknet_leaf_13_clk _0872_ VGND VGND VPWR VPWR rf.registers\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8514__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7639_ net151 _3464_ _3772_ VGND VGND VPWR VPWR _3777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7009__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9309_ clknet_leaf_14_clk _0469_ VGND VGND VPWR VPWR rf.registers\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6149__A _1731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7679__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7005__A1 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5111__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5319__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold109 rf.registers\[18\]\[18\] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4542__A2 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6758__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5178__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6059__A _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6493__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7990_ _3962_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6941_ _3390_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5350__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6872_ net214 _3118_ _3351_ VGND VGND VPWR VPWR _3354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8611_ clknet_leaf_68_clk _0795_ VGND VGND VPWR VPWR rf.registers\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5823_ _2472_ _2570_ _2571_ _1111_ VGND VGND VPWR VPWR _2572_ sky130_fd_sc_hd__a22o_1
X_9591_ clknet_leaf_26_clk _0751_ VGND VGND VPWR VPWR rf.registers\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8542_ _4254_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8213__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5754_ _1125_ _1110_ _1144_ _1166_ VGND VGND VPWR VPWR _2506_ sky130_fd_sc_hd__and4_1
XFILLER_0_134_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4705_ rf.registers\[12\]\[12\] rf.registers\[13\]\[12\] rf.registers\[14\]\[12\]
+ rf.registers\[15\]\[12\] net1155 _1183_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__mux4_1
X_8473_ net414 net17 _4216_ VGND VGND VPWR VPWR _4219_ sky130_fd_sc_hd__mux2_1
X_5685_ _2178_ _1802_ _2438_ VGND VGND VPWR VPWR _2439_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_20_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5138__A _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7424_ _3662_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__clkbuf_1
X_4636_ _1048_ _1391_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold610 rf.registers\[1\]\[14\] VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold621 rf.registers\[12\]\[2\] VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4977__A _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7355_ _3625_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_116_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4567_ _1319_ _1322_ _1213_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_116_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5572__S _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold632 rf.registers\[2\]\[20\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 rf.registers\[11\]\[17\] VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _3019_ net680 _3023_ VGND VGND VPWR VPWR _3024_ sky130_fd_sc_hd__mux2_1
Xhold654 rf.registers\[2\]\[30\] VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold665 rf.registers\[25\]\[8\] VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__dlygate4sd3_1
X_7286_ _3087_ net1061 _3554_ VGND VGND VPWR VPWR _3589_ sky130_fd_sc_hd__mux2_1
Xhold676 rf.registers\[8\]\[20\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _1205_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__buf_4
Xhold687 rf.registers\[25\]\[19\] VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd3_1
X_9025_ clknet_leaf_58_clk _0185_ VGND VGND VPWR VPWR rf.registers\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold698 rf.registers\[25\]\[27\] VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd3_1
X_6237_ _2701_ _2797_ VGND VGND VPWR VPWR _2964_ sky130_fd_sc_hd__nor2_1
X_6168_ _2390_ _2864_ _2333_ VGND VGND VPWR VPWR _2899_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7499__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5119_ _1758_ _1874_ _1800_ VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__o21ai_1
X_6099_ _2806_ _2827_ _2831_ _2833_ VGND VGND VPWR VPWR _2834_ sky130_fd_sc_hd__o31a_1
XANTENNA__5797__A1 _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8809_ clknet_leaf_47_clk _0993_ VGND VGND VPWR VPWR rf.registers\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone21 net108 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4772__A2 _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5990__B _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6578__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7263__A _3554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5688__B_N _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7202__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5332__S0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4460__B2 _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6342__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8033__S _3951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5960__A1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7872__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5470_ rf.registers\[0\]\[8\] rf.registers\[1\]\[8\] rf.registers\[2\]\[8\] rf.registers\[3\]\[8\]
+ _1734_ _1735_ VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4421_ rf.registers\[16\]\[29\] rf.registers\[17\]\[29\] rf.registers\[18\]\[29\]
+ rf.registers\[19\]\[29\] _1173_ _1175_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__mux4_2
XANTENNA__4797__A _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5712__A1 _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7140_ net241 _3444_ _3498_ VGND VGND VPWR VPWR _3511_ sky130_fd_sc_hd__mux2_1
X_4352_ _1103_ _1106_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7071_ net528 _3464_ _3456_ VGND VGND VPWR VPWR _3465_ sky130_fd_sc_hd__mux2_1
X_4283_ _1030_ _1031_ _1032_ _1033_ _1036_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__mux4_2
X_6022_ _1512_ _1587_ _2658_ _2741_ VGND VGND VPWR VPWR _2761_ sky130_fd_sc_hd__a31o_1
XANTENNA__4374__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4736__S _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7973_ _3095_ net1101 _3952_ VGND VGND VPWR VPWR _3954_ sky130_fd_sc_hd__mux2_1
X_6924_ _3381_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6855_ net708 _3101_ _3340_ VGND VGND VPWR VPWR _3345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4471__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5806_ _2496_ _2549_ _2552_ _2555_ VGND VGND VPWR VPWR _2556_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9574_ clknet_leaf_1_clk _0734_ VGND VGND VPWR VPWR rf.registers\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6786_ _3308_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8525_ net449 net41 _4244_ VGND VGND VPWR VPWR _4246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5737_ _1666_ _2488_ VGND VGND VPWR VPWR _2489_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8456_ net900 net40 _4205_ VGND VGND VPWR VPWR _4210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5668_ _1128_ _2420_ _2421_ VGND VGND VPWR VPWR _2422_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7407_ _3071_ rf.registers\[26\]\[23\] _3650_ VGND VGND VPWR VPWR _3654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4619_ _1371_ _1372_ _1373_ _1374_ _1190_ _1254_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__mux4_1
XANTENNA__6398__S _3022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8387_ _4173_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5599_ _2352_ _2353_ VGND VGND VPWR VPWR _2354_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold440 rf.registers\[25\]\[30\] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
X_7338_ _3071_ net262 _3613_ VGND VGND VPWR VPWR _3617_ sky130_fd_sc_hd__mux2_1
Xhold451 rf.registers\[10\]\[23\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 rf.registers\[0\]\[7\] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 rf.registers\[7\]\[7\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 rf.registers\[0\]\[30\] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold495 rf.registers\[7\]\[18\] VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
X_7269_ _3580_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9008_ clknet_leaf_3_clk _0168_ VGND VGND VPWR VPWR rf.registers\[31\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4365__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4646__S _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8118__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4690__A1 _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7957__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6861__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5477__S _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7392__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload18 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload29 clknet_leaf_57_clk VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_8
XFILLER_0_121_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4356__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5553__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output57_A net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5241__A _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4970_ _1685_ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5895__B _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6640_ _3003_ _3155_ VGND VGND VPWR VPWR _3230_ sky130_fd_sc_hd__nor2_4
XFILLER_0_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6571_ net10 net9 net46 VGND VGND VPWR VPWR _3193_ sky130_fd_sc_hd__and3_4
XFILLER_0_116_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8310_ _3090_ _3155_ VGND VGND VPWR VPWR _4132_ sky130_fd_sc_hd__nor2_4
XFILLER_0_82_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5522_ rf.registers\[12\]\[7\] rf.registers\[13\]\[7\] rf.registers\[14\]\[7\] rf.registers\[15\]\[7\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2278_ sky130_fd_sc_hd__mux4_1
X_9290_ clknet_leaf_64_clk _0450_ VGND VGND VPWR VPWR rf.registers\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8241_ _4095_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__clkbuf_1
X_5453_ _1828_ _2208_ _1728_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4404_ _1158_ _1159_ _1047_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__mux2_1
X_8172_ net244 _3452_ _4024_ VGND VGND VPWR VPWR _4059_ sky130_fd_sc_hd__mux2_1
X_5384_ _1670_ _2131_ _2135_ _2139_ VGND VGND VPWR VPWR _2140_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7123_ net27 VGND VGND VPWR VPWR _3500_ sky130_fd_sc_hd__buf_2
X_4335_ rf.registers\[20\]\[3\] rf.registers\[21\]\[3\] rf.registers\[22\]\[3\] rf.registers\[23\]\[3\]
+ net102 _1090_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6946__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7054_ net281 _3452_ _3412_ VGND VGND VPWR VPWR _3453_ sky130_fd_sc_hd__mux2_1
XANTENNA__4347__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6005_ _2663_ _2689_ _2712_ _2725_ VGND VGND VPWR VPWR _2745_ sky130_fd_sc_hd__or4_4
XANTENNA__7777__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6681__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7956_ _3944_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6907_ net798 _3013_ _3362_ VGND VGND VPWR VPWR _3372_ sky130_fd_sc_hd__mux2_1
X_7887_ _3145_ net1093 _3902_ VGND VGND VPWR VPWR _3908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6838_ _3335_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9557_ clknet_leaf_32_clk _0717_ VGND VGND VPWR VPWR rf.registers\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6769_ _3298_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4283__S0 _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8508_ net242 net35 _4227_ VGND VGND VPWR VPWR _4237_ sky130_fd_sc_hd__mux2_1
XANTENNA__8401__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9488_ clknet_leaf_10_clk _0648_ VGND VGND VPWR VPWR rf.registers\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7677__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8439_ _4200_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5326__A _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7017__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4586__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold270 rf.registers\[13\]\[0\] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 rf.registers\[1\]\[12\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 rf.registers\[2\]\[16\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5535__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7687__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4405__A _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__A1 _2390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4274__S0 _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7668__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5679__B1 _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5236__A _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6766__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5526__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 A1[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
X_7810_ _3867_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__clkbuf_1
X_8790_ clknet_leaf_24_clk _0974_ VGND VGND VPWR VPWR rf.registers\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7741_ _3064_ net1046 _3830_ VGND VGND VPWR VPWR _3831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4953_ rf.registers\[8\]\[23\] rf.registers\[9\]\[23\] rf.registers\[10\]\[23\] rf.registers\[11\]\[23\]
+ _1705_ _1708_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__mux4_1
XANTENNA__4501__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4315__A _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7672_ _3771_ VGND VGND VPWR VPWR _3794_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4884_ net5 VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__inv_2
X_9411_ clknet_leaf_54_clk _0571_ VGND VGND VPWR VPWR rf.registers\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6623_ _3221_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5906__A1 _2650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9342_ clknet_leaf_72_clk _0502_ VGND VGND VPWR VPWR rf.registers\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6554_ net986 _3143_ _3179_ VGND VGND VPWR VPWR _3184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5505_ _2259_ _2260_ _2044_ VGND VGND VPWR VPWR _2261_ sky130_fd_sc_hd__mux2_1
X_9273_ clknet_leaf_20_clk _0433_ VGND VGND VPWR VPWR rf.registers\[23\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6485_ net531 _3145_ _3135_ VGND VGND VPWR VPWR _3146_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8224_ net305 _3504_ _4083_ VGND VGND VPWR VPWR _4087_ sky130_fd_sc_hd__mux2_1
X_5436_ _1828_ _2191_ _1728_ VGND VGND VPWR VPWR _2192_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8155_ _4050_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__clkbuf_1
X_5367_ _1671_ _2110_ _2122_ VGND VGND VPWR VPWR _2123_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_100_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7106_ _3488_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8084__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4318_ rf.registers\[8\]\[5\] rf.registers\[9\]\[5\] rf.registers\[10\]\[5\] rf.registers\[11\]\[5\]
+ net106 _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__mux4_1
XANTENNA__5517__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8086_ net471 _3502_ _4011_ VGND VGND VPWR VPWR _4014_ sky130_fd_sc_hd__mux2_1
X_5298_ rf.registers\[8\]\[3\] rf.registers\[9\]\[3\] rf.registers\[10\]\[3\] rf.registers\[11\]\[3\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2054_ sky130_fd_sc_hd__mux4_1
X_7037_ _3441_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_126_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4740__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7300__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8988_ clknet_leaf_12_clk _0148_ VGND VGND VPWR VPWR rf.registers\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_7939_ _3935_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7536__A _3699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8131__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5384__A1_N _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6586__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5508__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8306__S _4096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7586__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6615__A _3194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7210__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4495__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4798__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6270_ _2991_ _2994_ VGND VGND VPWR VPWR _2995_ sky130_fd_sc_hd__xnor2_2
X_5221_ _1766_ _1976_ _1672_ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5152_ _1906_ _1907_ _1745_ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7813__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5083_ net82 VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__buf_2
XANTENNA__4627__A1 _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5824__A0 _2470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8911_ clknet_leaf_28_clk _0071_ VGND VGND VPWR VPWR rf.registers\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8842_ clknet_leaf_7_clk _0002_ VGND VGND VPWR VPWR rf.registers\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8773_ clknet_leaf_52_clk _0957_ VGND VGND VPWR VPWR rf.registers\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5985_ _2140_ net1165 VGND VGND VPWR VPWR _2726_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7724_ _3048_ net218 _3819_ VGND VGND VPWR VPWR _3822_ sky130_fd_sc_hd__mux2_1
X_4936_ _1691_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__buf_4
XANTENNA__7329__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7655_ _3785_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_10 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4867_ rf.registers\[24\]\[18\] rf.registers\[25\]\[18\] rf.registers\[26\]\[18\]
+ rf.registers\[27\]\[18\] net109 _1202_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__mux4_1
XANTENNA_21 _3771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6606_ _3212_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7586_ _3046_ net636 _3747_ VGND VGND VPWR VPWR _3749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4798_ rf.registers\[4\]\[10\] rf.registers\[5\]\[10\] rf.registers\[6\]\[10\] rf.registers\[7\]\[10\]
+ net107 _1105_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9325_ clknet_leaf_41_clk _0485_ VGND VGND VPWR VPWR rf.registers\[21\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6537_ net1057 _3126_ _3168_ VGND VGND VPWR VPWR _3175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7790__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9256_ clknet_leaf_47_clk _0416_ VGND VGND VPWR VPWR rf.registers\[23\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6468_ net26 VGND VGND VPWR VPWR _3134_ sky130_fd_sc_hd__buf_2
XFILLER_0_30_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8207_ net381 _3487_ _4072_ VGND VGND VPWR VPWR _4078_ sky130_fd_sc_hd__mux2_1
X_5419_ _1670_ _2166_ _2170_ _2174_ VGND VGND VPWR VPWR _2175_ sky130_fd_sc_hd__a2bb2o_2
X_9187_ clknet_leaf_66_clk _0347_ VGND VGND VPWR VPWR rf.registers\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6399_ _3086_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8138_ _4041_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6068__B1 _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7804__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8069_ net1070 _3485_ _4000_ VGND VGND VPWR VPWR _4005_ sky130_fd_sc_hd__mux2_1
XANTENNA__4713__S1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8126__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7030__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4477__S0 _1182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7965__S _3915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6791__A1 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5594__A2 _2175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6543__A1 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4829__S _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4857__A1 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8048__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4704__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6345__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8220__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5770_ _2503_ _2520_ VGND VGND VPWR VPWR _2521_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4721_ rf.registers\[0\]\[13\] rf.registers\[1\]\[13\] rf.registers\[2\]\[13\] rf.registers\[3\]\[13\]
+ net1161 _1279_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5395__S net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7440_ _3671_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4652_ rf.registers\[8\]\[7\] rf.registers\[9\]\[7\] rf.registers\[10\]\[7\] rf.registers\[11\]\[7\]
+ net120 _1193_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput30 WD3[24] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7371_ _3035_ net1105 _3628_ VGND VGND VPWR VPWR _3635_ sky130_fd_sc_hd__mux2_1
Xinput41 WD3[5] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
X_4583_ _1335_ _1336_ _1337_ _1338_ _1189_ _1205_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__mux4_2
XANTENNA__4640__S0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold803 rf.registers\[12\]\[12\] VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd3_1
X_9110_ clknet_leaf_24_clk _0270_ VGND VGND VPWR VPWR rf.registers\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6322_ _3034_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__clkbuf_1
Xhold814 rf.registers\[6\]\[21\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 rf.registers\[28\]\[16\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold836 rf.registers\[31\]\[22\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold847 rf.registers\[23\]\[8\] VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold858 rf.registers\[14\]\[14\] VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__dlygate4sd3_1
X_9041_ clknet_leaf_40_clk _0201_ VGND VGND VPWR VPWR rf.registers\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold869 rf.registers\[30\]\[7\] VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlygate4sd3_1
X_6253_ _2255_ _2910_ _2978_ VGND VGND VPWR VPWR _2979_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5196__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5204_ _1839_ _1959_ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__nor2_1
XANTENNA__5844__A1_N _2038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6184_ _2408_ _2906_ _2907_ _2913_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__o22a_2
XANTENNA__6954__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5135_ rf.registers\[8\]\[31\] rf.registers\[9\]\[31\] rf.registers\[10\]\[31\] rf.registers\[11\]\[31\]
+ _1882_ _1884_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5066_ _1782_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_123_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8825_ clknet_leaf_20_clk _1009_ VGND VGND VPWR VPWR rf.registers\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7785__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5968_ net88 _1480_ _1464_ _2411_ VGND VGND VPWR VPWR _2710_ sky130_fd_sc_hd__a31o_1
X_8756_ clknet_leaf_30_clk _0940_ VGND VGND VPWR VPWR rf.registers\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7707_ _3031_ net1035 _3808_ VGND VGND VPWR VPWR _3813_ sky130_fd_sc_hd__mux2_1
X_4919_ _1674_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_101_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5899_ _2642_ _2643_ VGND VGND VPWR VPWR _2644_ sky130_fd_sc_hd__nand2_1
X_8687_ clknet_leaf_9_clk _0871_ VGND VGND VPWR VPWR rf.registers\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4503__A _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7638_ _3776_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7722__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6525__A1 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7569_ _3029_ net894 _3736_ VGND VGND VPWR VPWR _3740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4631__S0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9308_ clknet_leaf_16_clk _0468_ VGND VGND VPWR VPWR rf.registers\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4649__S _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9239_ clknet_leaf_22_clk _0399_ VGND VGND VPWR VPWR rf.registers\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5334__A _1645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8450__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7695__S _3771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5111__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4870__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6516__A1 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4413__A _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5178__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6774__S _3266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6940_ net169 _3118_ _3387_ VGND VGND VPWR VPWR _3390_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5350__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6871_ _3353_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__clkbuf_1
X_8610_ clknet_leaf_55_clk _0794_ VGND VGND VPWR VPWR rf.registers\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5822_ _2474_ _2469_ _1126_ VGND VGND VPWR VPWR _2571_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9590_ clknet_leaf_25_clk _0750_ VGND VGND VPWR VPWR rf.registers\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8541_ net187 net18 _4244_ VGND VGND VPWR VPWR _4254_ sky130_fd_sc_hd__mux2_1
X_5753_ _2496_ _2502_ _2504_ VGND VGND VPWR VPWR _2505_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4704_ rf.registers\[8\]\[12\] rf.registers\[9\]\[12\] rf.registers\[10\]\[12\] rf.registers\[11\]\[12\]
+ net1155 _1183_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__mux4_1
X_8472_ _4218_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5684_ _1841_ _2347_ VGND VGND VPWR VPWR _2438_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7423_ _3087_ net744 _3627_ VGND VGND VPWR VPWR _3662_ sky130_fd_sc_hd__mux2_1
X_4635_ rf.registers\[8\]\[6\] rf.registers\[9\]\[6\] rf.registers\[10\]\[6\] rf.registers\[11\]\[6\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7354_ _3087_ net382 _3590_ VGND VGND VPWR VPWR _3625_ sky130_fd_sc_hd__mux2_1
Xhold600 rf.registers\[14\]\[23\] VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 rf.registers\[30\]\[9\] VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _1320_ _1321_ _1198_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold622 rf.registers\[16\]\[14\] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold633 rf.registers\[19\]\[0\] VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6305_ _3022_ VGND VGND VPWR VPWR _3023_ sky130_fd_sc_hd__clkbuf_8
Xhold644 rf.registers\[13\]\[18\] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 rf.registers\[0\]\[29\] VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__dlygate4sd3_1
X_7285_ _3588_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__9493__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4497_ _1251_ _1252_ _1211_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__mux2_1
Xhold666 rf.registers\[14\]\[25\] VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 rf.registers\[23\]\[19\] VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__dlygate4sd3_1
X_9024_ clknet_leaf_68_clk _0184_ VGND VGND VPWR VPWR rf.registers\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold688 rf.registers\[17\]\[19\] VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 rf.registers\[27\]\[24\] VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd3_1
X_6236_ _1087_ _2960_ _2961_ _2962_ _1127_ VGND VGND VPWR VPWR _2963_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_139_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6684__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6167_ _2105_ _2754_ _2897_ _1087_ VGND VGND VPWR VPWR _2898_ sky130_fd_sc_hd__o211a_1
XANTENNA__8432__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5118_ _1777_ _1865_ _1869_ _1873_ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__o2bb2a_2
X_6098_ _2830_ _2832_ _2503_ VGND VGND VPWR VPWR _2833_ sky130_fd_sc_hd__o21a_1
X_5049_ rf.registers\[20\]\[18\] rf.registers\[21\]\[18\] rf.registers\[22\]\[18\]
+ rf.registers\[23\]\[18\] _1719_ _1722_ VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__mux4_1
XANTENNA__6994__A1 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8808_ clknet_leaf_63_clk _0992_ VGND VGND VPWR VPWR rf.registers\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8739_ clknet_leaf_67_clk _0923_ VGND VGND VPWR VPWR rf.registers\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone11 A2[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone22 _1172_ VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_152_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone44 _1026_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6859__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4379__S _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5332__S1 _1655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7719__A _3807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8314__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7162__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4420_ rf.registers\[20\]\[29\] rf.registers\[21\]\[29\] rf.registers\[22\]\[29\]
+ rf.registers\[23\]\[29\] _1173_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4351_ _1034_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7070_ net40 VGND VGND VPWR VPWR _3464_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4282_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6021_ _2757_ _2731_ _2758_ _2759_ VGND VGND VPWR VPWR _2760_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_3_3__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8285__A _4096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7972_ _3953_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6923_ net842 _3101_ _3376_ VGND VGND VPWR VPWR _3381_ sky130_fd_sc_hd__mux2_1
XANTENNA__8224__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6854_ _3344_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5087__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5805_ _1666_ _2554_ VGND VGND VPWR VPWR _2555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6785_ net204 _3099_ _3304_ VGND VGND VPWR VPWR _3308_ sky130_fd_sc_hd__mux2_1
X_9573_ clknet_leaf_61_clk _0733_ VGND VGND VPWR VPWR rf.registers\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5936__C1 _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5149__A _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4834__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8524_ _4245_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__clkbuf_1
X_5736_ _2040_ _2486_ _2487_ _1962_ VGND VGND VPWR VPWR _2488_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_118_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8455_ _4209_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__clkbuf_1
X_5667_ _2333_ VGND VGND VPWR VPWR _2421_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6679__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7406_ _3653_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4618_ rf.registers\[20\]\[24\] rf.registers\[21\]\[24\] rf.registers\[22\]\[24\]
+ rf.registers\[23\]\[24\] _1360_ _1361_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__mux4_1
X_8386_ net442 _3462_ _4169_ VGND VGND VPWR VPWR _4173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5598_ _1668_ _2247_ VGND VGND VPWR VPWR _2353_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold430 rf.registers\[29\]\[7\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
X_7337_ _3616_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
Xhold441 rf.registers\[1\]\[3\] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _1303_ _1304_ _1259_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_147_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold452 rf.registers\[31\]\[12\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 rf.registers\[5\]\[26\] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold474 rf.registers\[7\]\[23\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 rf.registers\[29\]\[0\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
X_7268_ _3069_ net1141 _3577_ VGND VGND VPWR VPWR _3580_ sky130_fd_sc_hd__mux2_1
Xhold496 rf.registers\[2\]\[19\] VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9007_ clknet_leaf_9_clk _0167_ VGND VGND VPWR VPWR rf.registers\[31\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6219_ _2105_ _2802_ _2946_ _1085_ VGND VGND VPWR VPWR _2947_ sky130_fd_sc_hd__o211a_1
X_7199_ _3542_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_51_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5612__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6967__A1 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5078__S0 _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7973__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5059__A _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4898__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7144__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload19 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_106_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5553__S1 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5241__B _1996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8044__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5069__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7883__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6570_ net13 net12 net11 VGND VGND VPWR VPWR _3192_ sky130_fd_sc_hd__and3b_2
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5521_ _2273_ _2274_ _2275_ _2276_ _1711_ _1716_ VGND VGND VPWR VPWR _2277_ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8240_ net148 _3452_ _4060_ VGND VGND VPWR VPWR _4095_ sky130_fd_sc_hd__mux2_1
X_5452_ _2206_ _2207_ _1738_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4403_ rf.registers\[12\]\[0\] rf.registers\[13\]\[0\] rf.registers\[14\]\[0\] rf.registers\[15\]\[0\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_10_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8171_ _4058_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5383_ _1828_ _2138_ _1728_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7122_ _3499_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_4334_ _1043_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7053_ net38 VGND VGND VPWR VPWR _3452_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6004_ _1874_ _2743_ VGND VGND VPWR VPWR _2744_ sky130_fd_sc_hd__xor2_1
X_7955_ net606 _3508_ _3938_ VGND VGND VPWR VPWR _3944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6906_ _3371_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__clkbuf_1
X_7886_ _3907_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6837_ net292 _3011_ _3326_ VGND VGND VPWR VPWR _3335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4807__S0 _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9556_ clknet_leaf_30_clk _0716_ VGND VGND VPWR VPWR rf.registers\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_rebuffer9_A _1348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6768_ _3081_ net724 _3289_ VGND VGND VPWR VPWR _3298_ sky130_fd_sc_hd__mux2_1
XANTENNA__4283__S1 _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8507_ _4236_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5719_ _2347_ _1169_ _1905_ VGND VGND VPWR VPWR _2472_ sky130_fd_sc_hd__and3_2
X_9487_ clknet_leaf_8_clk _0647_ VGND VGND VPWR VPWR rf.registers\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6699_ _3261_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4511__A _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8438_ net589 net34 _4191_ VGND VGND VPWR VPWR _4200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5232__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8369_ _4163_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__clkbuf_1
Xhold260 rf.registers\[9\]\[22\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8629__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold271 rf.registers\[12\]\[7\] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 rf.registers\[19\]\[13\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold293 rf.registers\[19\]\[2\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4657__S _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8129__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6438__A _3092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5535__S1 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5342__A _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6872__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5299__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4274__S1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7117__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7208__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4567__S _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6348__A net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5526__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5567__A1_N _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 A2[2] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_0_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7740_ _3807_ VGND VGND VPWR VPWR _3830_ sky130_fd_sc_hd__clkbuf_8
X_4952_ _1707_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4883_ _1638_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__buf_4
X_7671_ _3793_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
X_9410_ clknet_leaf_55_clk _0570_ VGND VGND VPWR VPWR rf.registers\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8502__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6622_ _3071_ net1027 _3217_ VGND VGND VPWR VPWR _3221_ sky130_fd_sc_hd__mux2_1
XANTENNA__5462__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9341_ clknet_leaf_15_clk _0501_ VGND VGND VPWR VPWR rf.registers\[21\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6553_ _3183_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7108__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5504_ rf.registers\[24\]\[6\] rf.registers\[25\]\[6\] rf.registers\[26\]\[6\] rf.registers\[27\]\[6\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2260_ sky130_fd_sc_hd__mux4_1
XANTENNA__5119__B1 _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9272_ clknet_leaf_26_clk _0432_ VGND VGND VPWR VPWR rf.registers\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6484_ net31 VGND VGND VPWR VPWR _3145_ sky130_fd_sc_hd__buf_2
XANTENNA__5214__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5435_ _2189_ _2190_ _1738_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__mux2_1
X_8223_ _4086_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6957__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5366_ _2112_ _2116_ _2121_ _1828_ _1728_ VGND VGND VPWR VPWR _2122_ sky130_fd_sc_hd__a221o_1
X_8154_ net1100 _3502_ _4047_ VGND VGND VPWR VPWR _4050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4317_ _1043_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__clkbuf_4
X_7105_ net968 _3487_ _3477_ VGND VGND VPWR VPWR _3488_ sky130_fd_sc_hd__mux2_1
X_8085_ _4013_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__clkbuf_1
X_5297_ _2052_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__6258__A _1923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5162__A _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5517__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7036_ net259 _3145_ _3435_ VGND VGND VPWR VPWR _3441_ sky130_fd_sc_hd__mux2_1
XANTENNA__7788__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6692__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8987_ clknet_leaf_35_clk _0147_ VGND VGND VPWR VPWR rf.registers\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7089__A _3455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4506__A _1219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7938_ net256 _3491_ _3927_ VGND VGND VPWR VPWR _3935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7869_ _3898_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9539_ clknet_leaf_67_clk _0699_ VGND VGND VPWR VPWR rf.registers\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7028__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4879__C _1634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5771__S _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5508__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5072__A _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4416__A _1072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4495__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8322__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5220_ _1974_ _1975_ _1745_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5151_ rf.registers\[16\]\[30\] rf.registers\[17\]\[30\] rf.registers\[18\]\[30\]
+ rf.registers\[19\]\[30\] _1895_ _1897_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7274__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5082_ _1671_ _1829_ _1833_ _1837_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__a2bb2o_2
X_8910_ clknet_leaf_29_clk _0070_ VGND VGND VPWR VPWR rf.registers\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7401__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8841_ clknet_leaf_47_clk _0001_ VGND VGND VPWR VPWR rf.registers\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6017__S _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8772_ clknet_leaf_52_clk _0956_ VGND VGND VPWR VPWR rf.registers\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5984_ _2123_ _2724_ VGND VGND VPWR VPWR _2725_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7723_ _3821_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__clkbuf_1
X_4935_ _1690_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_111_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8232__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_11 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7654_ net228 _3479_ _3783_ VGND VGND VPWR VPWR _3785_ sky130_fd_sc_hd__mux2_1
X_4866_ rf.registers\[28\]\[18\] rf.registers\[29\]\[18\] rf.registers\[30\]\[18\]
+ rf.registers\[31\]\[18\] net109 _1202_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__mux4_1
XANTENNA_22 _3843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6605_ _3054_ net1115 _3206_ VGND VGND VPWR VPWR _3212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4797_ _1038_ _1552_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7585_ _3748_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9324_ clknet_leaf_50_clk _0484_ VGND VGND VPWR VPWR rf.registers\[21\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6536_ _3174_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9255_ clknet_leaf_66_clk _0415_ VGND VGND VPWR VPWR rf.registers\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8468__A _4204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6467_ _3133_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8206_ _4077_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__clkbuf_1
X_5418_ _1828_ _2173_ _1728_ VGND VGND VPWR VPWR _2174_ sky130_fd_sc_hd__a21oi_1
X_9186_ clknet_leaf_59_clk _0346_ VGND VGND VPWR VPWR rf.registers\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6398_ _3085_ net1078 _3022_ VGND VGND VPWR VPWR _3086_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_120_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8137_ net324 _3485_ _4036_ VGND VGND VPWR VPWR _4041_ sky130_fd_sc_hd__mux2_1
X_5349_ _2104_ VGND VGND VPWR VPWR _2105_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8068_ _4004_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5276__C1 _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7019_ net514 _3128_ _3424_ VGND VGND VPWR VPWR _3432_ sky130_fd_sc_hd__mux2_1
XANTENNA__8407__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7311__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4477__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5426__S0 _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7981__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5067__A _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6597__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8052__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4720_ rf.registers\[4\]\[13\] rf.registers\[5\]\[13\] rf.registers\[6\]\[13\] rf.registers\[7\]\[13\]
+ net1161 _1279_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4651_ rf.registers\[12\]\[7\] rf.registers\[13\]\[7\] rf.registers\[14\]\[7\] rf.registers\[15\]\[7\]
+ net120 _1193_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7891__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput20 WD3[15] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
Xinput31 WD3[25] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
X_7370_ _3634_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
X_4582_ rf.registers\[20\]\[30\] rf.registers\[21\]\[30\] rf.registers\[22\]\[30\]
+ rf.registers\[23\]\[30\] _1267_ _1268_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__mux4_2
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 WD3[6] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
XFILLER_0_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6321_ _3033_ net376 _3023_ VGND VGND VPWR VPWR _3034_ sky130_fd_sc_hd__mux2_1
Xhold804 rf.registers\[26\]\[7\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4640__S1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold815 rf.registers\[28\]\[17\] VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 rf.registers\[29\]\[8\] VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold837 rf.registers\[19\]\[19\] VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 rf.registers\[16\]\[5\] VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9040_ clknet_leaf_3_clk _0200_ VGND VGND VPWR VPWR rf.registers\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6252_ _2104_ _2849_ _2977_ _1086_ VGND VGND VPWR VPWR _2978_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold859 rf.registers\[28\]\[19\] VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5203_ _1842_ _1958_ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6183_ _2504_ _2908_ _2912_ VGND VGND VPWR VPWR _2913_ sky130_fd_sc_hd__or3_1
X_5134_ _1885_ _1886_ _1887_ _1888_ _1889_ _1773_ VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__mux4_1
XANTENNA__7798__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5065_ _1758_ _1820_ VGND VGND VPWR VPWR _1821_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_123_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6470__A1 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4481__B1 _1236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8824_ clknet_leaf_27_clk _1008_ VGND VGND VPWR VPWR rf.registers\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8755_ clknet_leaf_33_clk _0939_ VGND VGND VPWR VPWR rf.registers\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5967_ _2550_ _2591_ _2708_ VGND VGND VPWR VPWR _2709_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_137_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4490__S _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7706_ _3812_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_43_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4918_ _1673_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_101_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8686_ clknet_leaf_29_clk _0870_ VGND VGND VPWR VPWR rf.registers\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_32_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
X_5898_ _2193_ _2640_ _2641_ VGND VGND VPWR VPWR _2643_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5408__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7637_ net925 _3462_ _3772_ VGND VGND VPWR VPWR _3776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4849_ _1603_ _1604_ _1178_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7568_ _3739_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4631__S1 _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9307_ clknet_leaf_34_clk _0467_ VGND VGND VPWR VPWR rf.registers\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_151_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6519_ _3165_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__clkbuf_1
X_7499_ _3027_ net879 _3700_ VGND VGND VPWR VPWR _3703_ sky130_fd_sc_hd__mux2_1
XANTENNA__7306__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9238_ clknet_leaf_25_clk _0398_ VGND VGND VPWR VPWR rf.registers\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4395__S0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9169_ clknet_leaf_42_clk _0329_ VGND VGND VPWR VPWR rf.registers\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8137__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6880__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7961__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4870__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5525__A _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7216__S _3516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7477__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7740__A _3807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5260__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6870_ net142 _3116_ _3351_ VGND VGND VPWR VPWR _3353_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_62_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7401__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5821_ net81 _2251_ VGND VGND VPWR VPWR _2570_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_85_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8540_ _4253_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4604__A _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5752_ _2503_ VGND VGND VPWR VPWR _2504_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_4703_ _1287_ _1458_ _1088_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8471_ net146 net16 _4216_ VGND VGND VPWR VPWR _4218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5683_ _2036_ _1757_ _2347_ VGND VGND VPWR VPWR _2437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7422_ _3661_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8510__S _4204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4634_ _1386_ _1387_ _1388_ _1389_ _1048_ _1088_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__mux4_2
XFILLER_0_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4565_ rf.registers\[24\]\[31\] rf.registers\[25\]\[31\] rf.registers\[26\]\[31\]
+ rf.registers\[27\]\[31\] _1200_ _1202_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__mux4_2
X_7353_ _3624_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
Xhold601 rf.registers\[0\]\[22\] VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold612 rf.registers\[4\]\[6\] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 rf.registers\[10\]\[18\] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6304_ _3020_ _3021_ VGND VGND VPWR VPWR _3022_ sky130_fd_sc_hd__nand2_4
Xhold634 rf.registers\[0\]\[10\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold645 rf.registers\[27\]\[15\] VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 rf.registers\[26\]\[4\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd3_1
X_7284_ _3085_ net786 _3554_ VGND VGND VPWR VPWR _3588_ sky130_fd_sc_hd__mux2_1
X_4496_ rf.registers\[0\]\[20\] rf.registers\[1\]\[20\] rf.registers\[2\]\[20\] rf.registers\[3\]\[20\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__mux4_1
Xhold667 rf.registers\[16\]\[24\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__dlygate4sd3_1
X_9023_ clknet_leaf_74_clk _0183_ VGND VGND VPWR VPWR rf.registers\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold678 rf.registers\[23\]\[17\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6965__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold689 rf.registers\[10\]\[4\] VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4377__S0 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6235_ _2102_ _2692_ VGND VGND VPWR VPWR _2962_ sky130_fd_sc_hd__nor2_1
X_6166_ _2255_ _2821_ _2896_ _2337_ VGND VGND VPWR VPWR _2897_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5117_ _1700_ _1872_ _1671_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__o21ai_1
X_6097_ _2806_ _2827_ VGND VGND VPWR VPWR _2832_ sky130_fd_sc_hd__nor2_1
X_5048_ _1757_ _1802_ _1803_ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__mux2_1
XANTENNA__9018__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7796__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8807_ clknet_leaf_2_clk _0991_ VGND VGND VPWR VPWR rf.registers\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5403__C1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6999_ _3421_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8738_ clknet_leaf_60_clk _0922_ VGND VGND VPWR VPWR rf.registers\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone12 A2[0] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_16
X_8669_ clknet_leaf_13_clk _0853_ VGND VGND VPWR VPWR rf.registers\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone45 _1219_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_16
XANTENNA__5706__B1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7036__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8120__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7934__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5945__B1 _2160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8330__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4350_ rf.registers\[0\]\[3\] rf.registers\[1\]\[3\] rf.registers\[2\]\[3\] rf.registers\[3\]\[3\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4281_ net7 VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__buf_4
XANTENNA__6785__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4359__S0 _1042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6020_ _2102_ _2406_ VGND VGND VPWR VPWR _2759_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_3_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7971_ _3089_ net1103 _3952_ VGND VGND VPWR VPWR _3953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6922_ _3380_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6853_ net310 _3099_ _3340_ VGND VGND VPWR VPWR _3344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5804_ _2442_ _2487_ _2553_ _2040_ VGND VGND VPWR VPWR _2554_ sky130_fd_sc_hd__o22a_1
XANTENNA__5087__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4334__A _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9572_ clknet_leaf_63_clk _0732_ VGND VGND VPWR VPWR rf.registers\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6784_ _3307_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8523_ net771 net40 _4244_ VGND VGND VPWR VPWR _4245_ sky130_fd_sc_hd__mux2_1
XANTENNA__5149__B _1904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4834__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5735_ net81 _2251_ VGND VGND VPWR VPWR _2487_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8240__S _4060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8454_ net300 net39 _4205_ VGND VGND VPWR VPWR _4209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5666_ _2363_ _2417_ _2419_ VGND VGND VPWR VPWR _2420_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7405_ _3069_ net882 _3650_ VGND VGND VPWR VPWR _3653_ sky130_fd_sc_hd__mux2_1
XANTENNA__4598__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6361__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4617_ rf.registers\[16\]\[24\] rf.registers\[17\]\[24\] rf.registers\[18\]\[24\]
+ rf.registers\[19\]\[24\] _1360_ _1361_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8385_ _4172_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5597_ _1839_ _2211_ VGND VGND VPWR VPWR _2352_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_131_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold420 rf.registers\[4\]\[29\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4911__A1 _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold431 rf.registers\[5\]\[16\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
X_7336_ _3069_ net918 _3613_ VGND VGND VPWR VPWR _3616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4548_ rf.registers\[24\]\[27\] rf.registers\[25\]\[27\] rf.registers\[26\]\[27\]
+ rf.registers\[27\]\[27\] _1262_ _1263_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold442 rf.registers\[27\]\[17\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 rf.registers\[4\]\[15\] VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold464 rf.registers\[21\]\[30\] VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 rf.registers\[12\]\[1\] VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 rf.registers\[28\]\[26\] VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
X_7267_ _3579_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
X_4479_ _1233_ _1234_ _1189_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__mux2_1
Xhold497 rf.registers\[8\]\[3\] VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
X_9006_ clknet_leaf_44_clk _0166_ VGND VGND VPWR VPWR rf.registers\[31\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6218_ _2255_ _2867_ _2945_ _2337_ VGND VGND VPWR VPWR _2946_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_5_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7198_ net910 _3502_ _3539_ VGND VGND VPWR VPWR _3542_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _1731_ _2853_ VGND VGND VPWR VPWR _2881_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7613__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8415__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5078__S1 _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clone24_A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8150__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8341__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6352__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4589__S0 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4761__S0 _1065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4419__A _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5949__S _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7080__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4513__S0 net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4853__S _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5069__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5520_ rf.registers\[20\]\[7\] rf.registers\[21\]\[7\] rf.registers\[22\]\[7\] rf.registers\[23\]\[7\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__mux4_1
XANTENNA__5167__A1_N _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5451_ rf.registers\[0\]\[10\] rf.registers\[1\]\[10\] rf.registers\[2\]\[10\] rf.registers\[3\]\[10\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4402_ rf.registers\[8\]\[0\] rf.registers\[9\]\[0\] rf.registers\[10\]\[0\] rf.registers\[11\]\[0\]
+ net107 _1105_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_97_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8170_ net380 _3450_ _4024_ VGND VGND VPWR VPWR _4058_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5382_ _2136_ _2137_ _1738_ VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7121_ net184 _3497_ _3498_ VGND VGND VPWR VPWR _3499_ sky130_fd_sc_hd__mux2_1
X_4333_ _1041_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__buf_12
XANTENNA__7843__A0 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7052_ _3451_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6003_ _1587_ _2742_ VGND VGND VPWR VPWR _2743_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4329__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4752__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4409__B1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7071__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4763__S _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7954_ _3943_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5621__A2 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6905_ net284 _3011_ _3362_ VGND VGND VPWR VPWR _3371_ sky130_fd_sc_hd__mux2_1
X_7885_ _3143_ net1016 _3902_ VGND VGND VPWR VPWR _3907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5909__B1 _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6836_ _3334_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4807__S1 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9555_ clknet_leaf_32_clk _0715_ VGND VGND VPWR VPWR rf.registers\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6767_ _3297_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8506_ net904 net34 _4227_ VGND VGND VPWR VPWR _4236_ sky130_fd_sc_hd__mux2_1
X_5718_ _2469_ _2470_ _2251_ VGND VGND VPWR VPWR _2471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9486_ clknet_leaf_41_clk _0646_ VGND VGND VPWR VPWR rf.registers\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6698_ net1059 _3009_ _3253_ VGND VGND VPWR VPWR _3261_ sky130_fd_sc_hd__mux2_1
X_8437_ _4199_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5649_ _2397_ _2403_ net87 VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5232__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8368_ net757 _3444_ _4155_ VGND VGND VPWR VPWR _4163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold250 rf.registers\[17\]\[22\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7319_ _3052_ net290 _3602_ VGND VGND VPWR VPWR _3607_ sky130_fd_sc_hd__mux2_1
Xhold261 rf.registers\[19\]\[22\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4991__S0 _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold272 rf.registers\[9\]\[20\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
X_8299_ _4126_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold283 rf.registers\[18\]\[19\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 rf.registers\[22\]\[5\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5342__B _2097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4743__S0 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5299__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8145__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8562__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5009__S _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6876__A1 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7224__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output62_A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4734__S0 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 A2[3] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8250__A0 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6800__A1 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4951_ _1706_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7670_ net578 _3495_ _3783_ VGND VGND VPWR VPWR _3793_ sky130_fd_sc_hd__mux2_1
X_4882_ _1637_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__buf_8
XANTENNA__5367__A1 _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6621_ _3220_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5462__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9340_ clknet_leaf_16_clk _0500_ VGND VGND VPWR VPWR rf.registers\[21\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6552_ net1096 _3141_ _3179_ VGND VGND VPWR VPWR _3183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5503_ rf.registers\[28\]\[6\] rf.registers\[29\]\[6\] rf.registers\[30\]\[6\] rf.registers\[31\]\[6\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9271_ clknet_leaf_33_clk _0431_ VGND VGND VPWR VPWR rf.registers\[23\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6483_ _3144_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7923__A _3915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5214__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8222_ net870 _3502_ _4083_ VGND VGND VPWR VPWR _4086_ sky130_fd_sc_hd__mux2_1
X_5434_ rf.registers\[0\]\[11\] rf.registers\[1\]\[11\] rf.registers\[2\]\[11\] rf.registers\[3\]\[11\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8153_ _4049_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5365_ _2119_ _2120_ _1738_ VGND VGND VPWR VPWR _2121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7104_ net20 VGND VGND VPWR VPWR _3487_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4316_ _1041_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__buf_12
XFILLER_0_10_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8084_ net1111 _3500_ _4011_ VGND VGND VPWR VPWR _4013_ sky130_fd_sc_hd__mux2_1
X_5296_ _1690_ VGND VGND VPWR VPWR _2052_ sky130_fd_sc_hd__buf_4
XANTENNA__6973__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7035_ _3440_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4725__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8986_ clknet_leaf_37_clk _0146_ VGND VGND VPWR VPWR rf.registers\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7937_ _3934_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5150__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7868_ _3126_ net991 _3891_ VGND VGND VPWR VPWR _3898_ sky130_fd_sc_hd__mux2_1
XANTENNA__8544__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6819_ _3325_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7799_ _3861_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9538_ clknet_leaf_60_clk _0698_ VGND VGND VPWR VPWR rf.registers\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9469_ clknet_leaf_15_clk _0629_ VGND VGND VPWR VPWR rf.registers\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_154_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4668__S _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7979__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4716__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8535__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6849__A1 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5150_ rf.registers\[20\]\[30\] rf.registers\[21\]\[30\] rf.registers\[22\]\[30\]
+ rf.registers\[23\]\[30\] _1895_ _1897_ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7889__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6793__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5081_ _1717_ _1836_ _1729_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5380__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7026__A1 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8840_ clknet_leaf_62_clk _0000_ VGND VGND VPWR VPWR rf.registers\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5037__B1 _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8771_ clknet_leaf_52_clk _0955_ VGND VGND VPWR VPWR rf.registers\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5132__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5983_ _1511_ _2723_ VGND VGND VPWR VPWR _2724_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7722_ _3046_ net819 _3819_ VGND VGND VPWR VPWR _3821_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4934_ _1642_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7653_ _3784_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4865_ _1619_ _1620_ _1259_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__mux2_1
XANTENNA_12 clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_23 _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6604_ _3211_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4342__A _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7584_ _3043_ net890 _3747_ VGND VGND VPWR VPWR _3748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4796_ _1550_ _1551_ _1047_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9323_ clknet_leaf_2_clk _0483_ VGND VGND VPWR VPWR rf.registers\[21\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6535_ net853 _3124_ _3168_ VGND VGND VPWR VPWR _3174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9254_ clknet_leaf_0_clk _0414_ VGND VGND VPWR VPWR rf.registers\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5199__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6466_ net770 _3132_ _3114_ VGND VGND VPWR VPWR _3133_ sky130_fd_sc_hd__mux2_1
X_8205_ net692 _3485_ _4072_ VGND VGND VPWR VPWR _4077_ sky130_fd_sc_hd__mux2_1
X_5417_ _2171_ _2172_ _1738_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9185_ clknet_leaf_58_clk _0345_ VGND VGND VPWR VPWR rf.registers\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6397_ net37 VGND VGND VPWR VPWR _3085_ sky130_fd_sc_hd__clkbuf_2
X_8136_ _4040_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__clkbuf_1
X_5348_ _1111_ VGND VGND VPWR VPWR _2104_ sky130_fd_sc_hd__clkbuf_4
X_8067_ net573 _3483_ _4000_ VGND VGND VPWR VPWR _4004_ sky130_fd_sc_hd__mux2_1
X_5279_ _1799_ _2034_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__and2_1
X_7018_ _3431_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7017__A1 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5112__S _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8969_ clknet_leaf_50_clk _0129_ VGND VGND VPWR VPWR rf.registers\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5348__A _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7039__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5426__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_rebuffer34_A _1542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6878__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5083__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5811__A _2286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4427__A _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5114__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__8333__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8508__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4650_ _1402_ _1405_ _1038_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__mux2_2
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 A3[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5742__A1 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput21 WD3[16] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
X_4581_ rf.registers\[16\]\[30\] rf.registers\[17\]\[30\] rf.registers\[18\]\[30\]
+ rf.registers\[19\]\[30\] _1267_ _1268_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__mux4_2
Xinput32 WD3[26] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput43 WD3[7] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XFILLER_0_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6320_ net41 VGND VGND VPWR VPWR _3033_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold805 rf.registers\[10\]\[25\] VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold816 rf.registers\[20\]\[11\] VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold827 rf.registers\[13\]\[22\] VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 rf.registers\[1\]\[10\] VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _1944_ _2975_ _2976_ VGND VGND VPWR VPWR _2977_ sky130_fd_sc_hd__o21ai_1
Xhold849 rf.registers\[6\]\[31\] VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5202_ _1777_ _1949_ _1957_ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__a21oi_2
X_6182_ _2530_ _2779_ _2911_ _1087_ VGND VGND VPWR VPWR _2912_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5133_ _1713_ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__buf_4
XANTENNA__8508__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5258__B1 _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5353__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5064_ _1671_ _1811_ _1815_ _1819_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_123_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4481__A1 _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5105__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8823_ clknet_leaf_24_clk _1007_ VGND VGND VPWR VPWR rf.registers\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8754_ clknet_leaf_28_clk _0938_ VGND VGND VPWR VPWR rf.registers\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5966_ _2553_ _2588_ _2679_ _2442_ _2333_ VGND VGND VPWR VPWR _2708_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7705_ _3029_ net1043 _3808_ VGND VGND VPWR VPWR _3812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4917_ _1641_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8685_ clknet_leaf_8_clk _0869_ VGND VGND VPWR VPWR rf.registers\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5897_ _2640_ _2641_ _2193_ VGND VGND VPWR VPWR _2642_ sky130_fd_sc_hd__a21o_1
XANTENNA__5981__B2 _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5168__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5408__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7636_ _3775_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_138_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4848_ rf.registers\[16\]\[19\] rf.registers\[17\]\[19\] rf.registers\[18\]\[19\]
+ rf.registers\[19\]\[19\] net127 _1222_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6698__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7567_ _3027_ net874 _3736_ VGND VGND VPWR VPWR _3739_ sky130_fd_sc_hd__mux2_1
X_4779_ _1047_ _1534_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__or2_4
XANTENNA__5733__B2 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9306_ clknet_leaf_37_clk _0466_ VGND VGND VPWR VPWR rf.registers\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6518_ net544 _3107_ _3157_ VGND VGND VPWR VPWR _3165_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7498_ _3702_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
X_9237_ clknet_leaf_31_clk _0397_ VGND VGND VPWR VPWR rf.registers\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6449_ _3121_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__clkbuf_1
X_9168_ clknet_leaf_12_clk _0328_ VGND VGND VPWR VPWR rf.registers\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4395__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8119_ _4031_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__clkbuf_1
X_9099_ clknet_leaf_3_clk _0259_ VGND VGND VPWR VPWR rf.registers\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5631__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6749__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5777__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4681__S _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6462__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7992__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5185__C1 _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6401__S _3022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5488__B1 _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8328__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7232__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5335__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5260__B _2015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7468__A _3663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8063__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5820_ _2568_ VGND VGND VPWR VPWR _2569_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5751_ net48 VGND VGND VPWR VPWR _2503_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_151_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4702_ rf.registers\[0\]\[12\] rf.registers\[1\]\[12\] rf.registers\[2\]\[12\] rf.registers\[3\]\[12\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__mux4_1
X_8470_ _4217_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__clkbuf_1
X_5682_ _2105_ _2427_ _2435_ VGND VGND VPWR VPWR _2436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7421_ _3085_ net1153 _3627_ VGND VGND VPWR VPWR _3661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4633_ rf.registers\[20\]\[6\] rf.registers\[21\]\[6\] rf.registers\[22\]\[6\] rf.registers\[23\]\[6\]
+ _1219_ _1221_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__mux4_2
XFILLER_0_154_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7407__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7352_ _3085_ net961 _3590_ VGND VGND VPWR VPWR _3624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4564_ rf.registers\[28\]\[31\] rf.registers\[29\]\[31\] rf.registers\[30\]\[31\]
+ rf.registers\[31\]\[31\] _1200_ _1202_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__mux4_1
Xhold602 rf.registers\[14\]\[8\] VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold613 rf.registers\[24\]\[16\] VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ net12 net11 net13 VGND VGND VPWR VPWR _3021_ sky130_fd_sc_hd__and3b_4
XTAP_TAPCELL_ROW_116_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold624 rf.registers\[3\]\[21\] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold635 rf.registers\[3\]\[9\] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__dlygate4sd3_1
X_7283_ _3587_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
Xhold646 rf.registers\[10\]\[0\] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ rf.registers\[4\]\[20\] rf.registers\[5\]\[20\] rf.registers\[6\]\[20\] rf.registers\[7\]\[20\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__mux4_1
Xhold657 rf.registers\[23\]\[14\] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlygate4sd3_1
X_9022_ clknet_leaf_74_clk _0182_ VGND VGND VPWR VPWR rf.registers\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold668 rf.registers\[31\]\[6\] VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 rf.registers\[24\]\[17\] VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _1111_ _2822_ _2896_ _2254_ VGND VGND VPWR VPWR _2961_ sky130_fd_sc_hd__o22a_1
XANTENNA__4377__S1 _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6165_ _2857_ _2895_ _2327_ VGND VGND VPWR VPWR _2896_ sky130_fd_sc_hd__mux2_1
XANTENNA__8238__S _4060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7142__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5116_ _1870_ _1871_ _1726_ VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__mux2_1
X_6096_ _2830_ VGND VGND VPWR VPWR _2831_ sky130_fd_sc_hd__inv_2
X_5047_ _1145_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5651__A0 _2390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8806_ clknet_leaf_2_clk _0990_ VGND VGND VPWR VPWR rf.registers\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6998_ net591 _3107_ _3413_ VGND VGND VPWR VPWR _3421_ sky130_fd_sc_hd__mux2_1
X_8737_ clknet_leaf_60_clk _0921_ VGND VGND VPWR VPWR rf.registers\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5949_ _2378_ _2381_ _2178_ VGND VGND VPWR VPWR _2692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8668_ clknet_leaf_18_clk _0852_ VGND VGND VPWR VPWR rf.registers\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xclone13 _1181_ VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__clkbuf_16
Xclone24 net108 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_16
Xclone35 net93 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone46 _1219_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_16
X_7619_ _3079_ net1098 _3758_ VGND VGND VPWR VPWR _3766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8599_ clknet_leaf_33_clk _0783_ VGND VGND VPWR VPWR rf.registers\[22\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7317__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5361__A _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7987__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6891__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6198__A1 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5300__S _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4280_ _1035_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__buf_6
XANTENNA__4359__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5556__S0 _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8058__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6367__A _3022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7897__S _3879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7970_ _3951_ VGND VGND VPWR VPWR _3952_ sky130_fd_sc_hd__clkbuf_8
X_6921_ net247 _3099_ _3376_ VGND VGND VPWR VPWR _3380_ sky130_fd_sc_hd__mux2_1
X_6852_ _3343_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6306__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5803_ _2443_ _2437_ _1879_ VGND VGND VPWR VPWR _2553_ sky130_fd_sc_hd__mux2_2
X_9571_ clknet_leaf_68_clk _0731_ VGND VGND VPWR VPWR rf.registers\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6783_ net378 _3097_ _3304_ VGND VGND VPWR VPWR _3307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8522_ _3006_ VGND VGND VPWR VPWR _4244_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5734_ _2037_ _1804_ _2251_ VGND VGND VPWR VPWR _2486_ sky130_fd_sc_hd__mux2_2
XFILLER_0_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7689__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8453_ _4208_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__clkbuf_1
X_5665_ _1147_ _2418_ VGND VGND VPWR VPWR _2419_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7404_ _3652_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__clkbuf_1
X_4616_ rf.registers\[28\]\[24\] rf.registers\[29\]\[24\] rf.registers\[30\]\[24\]
+ rf.registers\[31\]\[24\] _1360_ _1361_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__mux4_1
X_8384_ net703 _3460_ _4169_ VGND VGND VPWR VPWR _4172_ sky130_fd_sc_hd__mux2_1
XANTENNA__4598__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5596_ _2349_ _2350_ VGND VGND VPWR VPWR _2351_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold410 rf.registers\[15\]\[26\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7335_ _3615_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
Xhold421 rf.registers\[26\]\[14\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ rf.registers\[28\]\[27\] rf.registers\[29\]\[27\] rf.registers\[30\]\[27\]
+ rf.registers\[31\]\[27\] _1262_ _1263_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__mux4_2
Xhold432 rf.registers\[19\]\[17\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 rf.registers\[1\]\[29\] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold454 rf.registers\[11\]\[21\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7266_ _3067_ net1138 _3577_ VGND VGND VPWR VPWR _3579_ sky130_fd_sc_hd__mux2_1
Xhold465 rf.registers\[24\]\[29\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 rf.registers\[0\]\[11\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ rf.registers\[12\]\[28\] rf.registers\[13\]\[28\] rf.registers\[14\]\[28\]
+ rf.registers\[15\]\[28\] _1182_ _1184_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__mux4_1
Xhold487 rf.registers\[9\]\[7\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9005_ clknet_leaf_41_clk _0165_ VGND VGND VPWR VPWR rf.registers\[31\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold498 rf.registers\[21\]\[16\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
X_6217_ _2909_ _2944_ _2178_ VGND VGND VPWR VPWR _2945_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7197_ _3541_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_51_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _1731_ _2853_ _2838_ VGND VGND VPWR VPWR _2880_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_51_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _2667_ net124 VGND VGND VPWR VPWR _2815_ sky130_fd_sc_hd__or2_1
XANTENNA__7600__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5356__A _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4589__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4559__A1_N _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6886__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_61_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5538__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6187__A _1978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4761__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4513__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4435__A _1072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6126__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4277__S0 _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__8341__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5450_ rf.registers\[4\]\[10\] rf.registers\[5\]\[10\] rf.registers\[6\]\[10\] rf.registers\[7\]\[10\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4401_ _1038_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5381_ rf.registers\[0\]\[14\] rf.registers\[1\]\[14\] rf.registers\[2\]\[14\] rf.registers\[3\]\[14\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2137_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_97_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7120_ _3455_ VGND VGND VPWR VPWR _3498_ sky130_fd_sc_hd__buf_4
X_4332_ _1050_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7051_ net393 _3450_ _3412_ VGND VGND VPWR VPWR _3451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6002_ _1512_ _2658_ _2741_ VGND VGND VPWR VPWR _2742_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4752__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8516__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4409__A1 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7953_ net942 _3506_ _3938_ VGND VGND VPWR VPWR _3943_ sky130_fd_sc_hd__mux2_1
X_6904_ _3370_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__clkbuf_1
X_7884_ _3906_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6835_ net351 _3009_ _3326_ VGND VGND VPWR VPWR _3334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9554_ clknet_leaf_27_clk _0714_ VGND VGND VPWR VPWR rf.registers\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6766_ _3079_ net700 _3289_ VGND VGND VPWR VPWR _3297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4999__B _1754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5717_ _2396_ _2400_ _1877_ VGND VGND VPWR VPWR _2470_ sky130_fd_sc_hd__mux2_1
X_8505_ _4235_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__clkbuf_1
X_9485_ clknet_leaf_40_clk _0645_ VGND VGND VPWR VPWR rf.registers\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6697_ _3260_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__clkbuf_1
X_5648_ _2400_ _2402_ _1145_ VGND VGND VPWR VPWR _2403_ sky130_fd_sc_hd__mux2_1
X_8436_ net576 net33 _4191_ VGND VGND VPWR VPWR _4199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8367_ _4162_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__clkbuf_1
X_5579_ _1128_ _1663_ _2334_ _2330_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__o211ai_4
XANTENNA__4440__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7318_ _3606_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
Xhold240 rf.registers\[22\]\[17\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold251 rf.registers\[9\]\[1\] VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 rf.registers\[10\]\[8\] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
X_8298_ _3002_ net1087 _4119_ VGND VGND VPWR VPWR _4126_ sky130_fd_sc_hd__mux2_1
Xhold273 rf.registers\[11\]\[10\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4991__S1 _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6098__B1 _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold284 rf.registers\[24\]\[5\] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 rf.registers\[26\]\[8\] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
X_7249_ _3050_ net504 _3566_ VGND VGND VPWR VPWR _3570_ sky130_fd_sc_hd__mux2_1
XANTENNA__4743__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8426__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8675__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5086__A _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7505__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7825__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4734__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 A2[4] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_4
XANTENNA__7240__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4950_ _1678_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4881_ _1448_ _1350_ _1385_ _1636_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__or4b_4
XFILLER_0_52_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6620_ _3069_ net884 _3217_ VGND VGND VPWR VPWR _3220_ sky130_fd_sc_hd__mux2_1
XANTENNA__8071__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6564__A1 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6551_ _3182_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5935__C_N _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5502_ _2256_ _2257_ _2044_ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4670__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9270_ clknet_leaf_24_clk _0430_ VGND VGND VPWR VPWR rf.registers\[23\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5119__A2 _1874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6482_ net509 _3143_ _3135_ VGND VGND VPWR VPWR _3144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8221_ _4085_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__clkbuf_1
X_5433_ rf.registers\[4\]\[11\] rf.registers\[5\]\[11\] rf.registers\[6\]\[11\] rf.registers\[7\]\[11\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2189_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7415__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8069__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8152_ net845 _3500_ _4047_ VGND VGND VPWR VPWR _4049_ sky130_fd_sc_hd__mux2_1
X_5364_ rf.registers\[0\]\[15\] rf.registers\[1\]\[15\] rf.registers\[2\]\[15\] rf.registers\[3\]\[15\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7103_ _3486_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_4315_ _1037_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8083_ _4012_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__clkbuf_1
X_5295_ _2050_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__buf_4
X_7034_ net285 _3143_ _3435_ VGND VGND VPWR VPWR _3440_ sky130_fd_sc_hd__mux2_1
XANTENNA__4725__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8246__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8985_ clknet_leaf_19_clk _0145_ VGND VGND VPWR VPWR rf.registers\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_7936_ net196 _3489_ _3927_ VGND VGND VPWR VPWR _3934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5150__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7867_ _3897_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6818_ net766 _3132_ _3315_ VGND VGND VPWR VPWR _3325_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7798_ net810 _3487_ _3855_ VGND VGND VPWR VPWR _3861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9537_ clknet_leaf_61_clk _0697_ VGND VGND VPWR VPWR rf.registers\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4522__B _1277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6749_ _3062_ net1125 _3278_ VGND VGND VPWR VPWR _3288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4661__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9468_ clknet_leaf_16_clk _0628_ VGND VGND VPWR VPWR rf.registers\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8419_ net466 _3495_ _4180_ VGND VGND VPWR VPWR _4190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7325__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9399_ clknet_leaf_34_clk _0559_ VGND VGND VPWR VPWR rf.registers\[24\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4716__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8156__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6465__A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6546__A1 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4652__S0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5544__A _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8471__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5080_ _1834_ _1835_ _1686_ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__mux2_1
XANTENNA__5285__A1 _2038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5380__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5037__A1 _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6785__A1 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8770_ clknet_leaf_55_clk _0954_ VGND VGND VPWR VPWR rf.registers\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_5982_ _1495_ net89 _2536_ VGND VGND VPWR VPWR _2723_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5132__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7721_ _3820_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__clkbuf_1
X_4933_ _1675_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_121_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4891__S0 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4623__A _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7652_ net361 _3476_ _3783_ VGND VGND VPWR VPWR _3784_ sky130_fd_sc_hd__mux2_1
X_4864_ rf.registers\[16\]\[18\] rf.registers\[17\]\[18\] rf.registers\[18\]\[18\]
+ rf.registers\[19\]\[18\] net109 _1202_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__mux4_1
XANTENNA__6537__A1 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_24 _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _3052_ net783 _3206_ VGND VGND VPWR VPWR _3211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7583_ _3735_ VGND VGND VPWR VPWR _3747_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4795_ rf.registers\[12\]\[10\] rf.registers\[13\]\[10\] rf.registers\[14\]\[10\]
+ rf.registers\[15\]\[10\] net117 _1090_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9322_ clknet_leaf_64_clk _0482_ VGND VGND VPWR VPWR rf.registers\[21\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6534_ _3173_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9253_ clknet_leaf_62_clk _0413_ VGND VGND VPWR VPWR rf.registers\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6465_ net24 VGND VGND VPWR VPWR _3132_ sky130_fd_sc_hd__buf_2
XANTENNA__5199__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5416_ rf.registers\[0\]\[12\] rf.registers\[1\]\[12\] rf.registers\[2\]\[12\] rf.registers\[3\]\[12\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__mux4_1
X_8204_ _4076_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__clkbuf_1
X_9184_ clknet_leaf_60_clk _0344_ VGND VGND VPWR VPWR rf.registers\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6396_ _3084_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8135_ net166 _3483_ _4036_ VGND VGND VPWR VPWR _4040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6984__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5347_ _1127_ _1663_ _2100_ _2102_ VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__a31o_1
XANTENNA__8462__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8066_ _4003_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__clkbuf_1
X_5278_ _1639_ _2033_ VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_34_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5276__B2 _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7017_ net1129 _3126_ _3424_ VGND VGND VPWR VPWR _3431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7973__A0 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8968_ clknet_leaf_46_clk _0128_ VGND VGND VPWR VPWR rf.registers\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_7919_ net401 _3472_ _3916_ VGND VGND VPWR VPWR _3925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8899_ clknet_leaf_52_clk _0059_ VGND VGND VPWR VPWR rf.registers\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5629__A _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4533__A _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4634__S0 _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6700__A1 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9219__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8205__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5114__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4443__A _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4625__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput11 A3[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4580_ rf.registers\[28\]\[30\] rf.registers\[29\]\[30\] rf.registers\[30\]\[30\]
+ rf.registers\[31\]\[30\] _1201_ _1203_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__mux4_2
Xinput22 WD3[17] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput33 WD3[27] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
Xinput44 WD3[8] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold806 rf.registers\[27\]\[31\] VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold817 rf.registers\[25\]\[21\] VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold828 rf.registers\[7\]\[22\] VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6250_ _2178_ _1980_ _1960_ _1127_ VGND VGND VPWR VPWR _2976_ sky130_fd_sc_hd__o31a_1
Xhold839 rf.registers\[14\]\[30\] VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5050__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5201_ _1951_ _1953_ _1956_ _1773_ _1672_ VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__o221a_2
XFILLER_0_110_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6181_ _2254_ _2848_ _2910_ _2336_ VGND VGND VPWR VPWR _2911_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5132_ rf.registers\[20\]\[31\] rf.registers\[21\]\[31\] rf.registers\[22\]\[31\]
+ rf.registers\[23\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__mux4_1
XANTENNA__8444__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5258__A1 _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6309__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5063_ _1717_ _1818_ _1729_ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5213__S _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5353__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8822_ clknet_leaf_24_clk _1006_ VGND VGND VPWR VPWR rf.registers\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5105__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5966__C1 _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8753_ clknet_leaf_29_clk _0937_ VGND VGND VPWR VPWR rf.registers\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5965_ _1087_ _2706_ VGND VGND VPWR VPWR _2707_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5449__A _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7704_ _3811_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4916_ _1671_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__buf_4
X_5896_ _2595_ _2639_ _1572_ VGND VGND VPWR VPWR _2641_ sky130_fd_sc_hd__a21o_1
X_8684_ clknet_leaf_63_clk _0868_ VGND VGND VPWR VPWR rf.registers\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5168__B _1923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7635_ net392 _3460_ _3772_ VGND VGND VPWR VPWR _3775_ sky130_fd_sc_hd__mux2_1
XANTENNA__6979__S _3375_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7183__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4847_ rf.registers\[20\]\[19\] rf.registers\[21\]\[19\] rf.registers\[22\]\[19\]
+ rf.registers\[23\]\[19\] net135 _1184_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7566_ _3738_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
X_4778_ rf.registers\[8\]\[9\] rf.registers\[9\]\[9\] rf.registers\[10\]\[9\] rf.registers\[11\]\[9\]
+ net107 _1105_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__mux4_2
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9305_ clknet_leaf_20_clk _0465_ VGND VGND VPWR VPWR rf.registers\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6517_ _3164_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_151_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7497_ _3025_ net676 _3700_ VGND VGND VPWR VPWR _3702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9236_ clknet_leaf_30_clk _0396_ VGND VGND VPWR VPWR rf.registers\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6448_ net415 _3120_ _3114_ VGND VGND VPWR VPWR _3121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9167_ clknet_leaf_28_clk _0327_ VGND VGND VPWR VPWR rf.registers\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6379_ net30 VGND VGND VPWR VPWR _3073_ sky130_fd_sc_hd__clkbuf_2
X_8118_ net366 _3466_ _4025_ VGND VGND VPWR VPWR _4031_ sky130_fd_sc_hd__mux2_1
X_9098_ clknet_leaf_8_clk _0258_ VGND VGND VPWR VPWR rf.registers\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8049_ _3994_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8434__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6889__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6921__A1 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5488__A1 _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_60_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7513__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8426__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4438__A _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5335__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5033__S _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__S _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5099__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5750_ _2497_ _2500_ _2501_ VGND VGND VPWR VPWR _2502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4701_ _1198_ _1456_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5681_ _2255_ _2431_ _2434_ _2373_ VGND VGND VPWR VPWR _2435_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4632_ rf.registers\[16\]\[6\] rf.registers\[17\]\[6\] rf.registers\[18\]\[6\] rf.registers\[19\]\[6\]
+ _1219_ _1221_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__mux4_2
XFILLER_0_72_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7420_ _3660_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5271__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4563_ _1317_ _1318_ _1198_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__mux2_1
X_7351_ _3623_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold603 rf.registers\[17\]\[11\] VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6302_ net9 _3004_ VGND VGND VPWR VPWR _3020_ sky130_fd_sc_hd__nor2_4
Xhold614 rf.registers\[20\]\[23\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold625 rf.registers\[13\]\[1\] VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7282_ _3083_ net912 _3577_ VGND VGND VPWR VPWR _3587_ sky130_fd_sc_hd__mux2_1
Xhold636 rf.registers\[28\]\[30\] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _1199_ _1249_ _1213_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold647 rf.registers\[14\]\[6\] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 rf.registers\[9\]\[21\] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9021_ clknet_leaf_3_clk _0181_ VGND VGND VPWR VPWR rf.registers\[31\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6233_ _1148_ _2958_ _2959_ _2337_ VGND VGND VPWR VPWR _2960_ sky130_fd_sc_hd__a211o_1
Xhold669 rf.registers\[31\]\[15\] VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7423__S _3627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8417__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6164_ _2386_ _2391_ VGND VGND VPWR VPWR _2895_ sky130_fd_sc_hd__nor2_1
X_5115_ rf.registers\[0\]\[16\] rf.registers\[1\]\[16\] rf.registers\[2\]\[16\] rf.registers\[3\]\[16\]
+ _1822_ _1823_ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__mux4_1
XANTENNA__4348__A _1041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6095_ _1779_ _2829_ VGND VGND VPWR VPWR _2830_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5046_ _1781_ _1801_ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_108_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8254__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8805_ clknet_leaf_53_clk _0989_ VGND VGND VPWR VPWR rf.registers\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6997_ _3420_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5179__A _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5403__B2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4837__S0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8736_ clknet_leaf_70_clk _0920_ VGND VGND VPWR VPWR rf.registers\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_5948_ _2661_ _2669_ _2689_ VGND VGND VPWR VPWR _2691_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8667_ clknet_leaf_23_clk _0851_ VGND VGND VPWR VPWR rf.registers\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5879_ _2548_ _2624_ _2426_ VGND VGND VPWR VPWR _2625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone25 net108 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_16
XANTENNA__4811__A _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7618_ _3765_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5706__A2 _2458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8598_ clknet_leaf_24_clk _0782_ VGND VGND VPWR VPWR rf.registers\[22\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5262__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7549_ _3077_ net1104 _3722_ VGND VGND VPWR VPWR _3729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5014__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9219_ clknet_leaf_68_clk _0379_ VGND VGND VPWR VPWR rf.registers\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8164__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4828__S0 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_135_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8339__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5556__S1 _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7243__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6920_ _3379_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6851_ net222 _3097_ _3340_ VGND VGND VPWR VPWR _3343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4819__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5802_ _2530_ _2550_ _2551_ _2373_ VGND VGND VPWR VPWR _2552_ sky130_fd_sc_hd__o211a_1
X_9570_ clknet_leaf_60_clk _0730_ VGND VGND VPWR VPWR rf.registers\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6782_ _3306_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8521_ _4243_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5733_ _2459_ _2467_ _2477_ _2485_ _2408_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__o32a_2
XFILLER_0_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5727__A _2062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8452_ net499 net36 _4205_ VGND VGND VPWR VPWR _4208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5664_ _2082_ _2099_ VGND VGND VPWR VPWR _2418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5244__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7403_ _3067_ net1119 _3650_ VGND VGND VPWR VPWR _3652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4615_ rf.registers\[24\]\[24\] rf.registers\[25\]\[24\] rf.registers\[26\]\[24\]
+ rf.registers\[27\]\[24\] _1360_ _1361_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8383_ _4171_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__clkbuf_1
X_5595_ _1668_ _2194_ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold400 rf.registers\[18\]\[14\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold411 rf.registers\[29\]\[4\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
X_7334_ _3067_ net877 _3613_ VGND VGND VPWR VPWR _3615_ sky130_fd_sc_hd__mux2_1
X_4546_ _1300_ _1301_ _1259_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__mux2_1
Xhold422 rf.registers\[29\]\[13\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 rf.registers\[11\]\[6\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 rf.registers\[20\]\[5\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 rf.registers\[20\]\[7\] VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 rf.registers\[26\]\[16\] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
X_7265_ _3578_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
X_4477_ rf.registers\[8\]\[28\] rf.registers\[9\]\[28\] rf.registers\[10\]\[28\] rf.registers\[11\]\[28\]
+ _1182_ _1184_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__mux4_1
Xhold477 rf.registers\[19\]\[9\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
X_9004_ clknet_leaf_49_clk _0164_ VGND VGND VPWR VPWR rf.registers\[31\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold488 rf.registers\[8\]\[14\] VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 rf.registers\[20\]\[10\] VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__dlygate4sd3_1
X_6216_ _1980_ _1960_ VGND VGND VPWR VPWR _2944_ sky130_fd_sc_hd__nor2_1
X_7196_ net911 _3500_ _3539_ VGND VGND VPWR VPWR _3541_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6992__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6147_ _2814_ _2815_ _2748_ _2816_ _2878_ VGND VGND VPWR VPWR _2879_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_51_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _2813_ _2665_ _2745_ _2600_ VGND VGND VPWR VPWR _2814_ sky130_fd_sc_hd__or4b_4
X_5029_ _1783_ _1784_ _1739_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5483__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8719_ clknet_leaf_28_clk _0903_ VGND VGND VPWR VPWR rf.registers\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5637__A _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5235__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6468__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5538__S1 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7998__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5311__S _1645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4277__S1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7238__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4451__A _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5226__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4400_ _1154_ _1155_ _1107_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4354__A1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5380_ rf.registers\[4\]\[14\] rf.registers\[5\]\[14\] rf.registers\[6\]\[14\] rf.registers\[7\]\[14\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_97_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4331_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__8069__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7050_ net37 VGND VGND VPWR VPWR _3450_ sky130_fd_sc_hd__buf_2
XFILLER_0_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6001_ _2536_ VGND VGND VPWR VPWR _2741_ sky130_fd_sc_hd__buf_2
XANTENNA__7701__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7952_ _3942_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6903_ net307 _3009_ _3362_ VGND VGND VPWR VPWR _3370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7883_ _3141_ net767 _3902_ VGND VGND VPWR VPWR _3906_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6834_ _3333_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5909__A2 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5465__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9553_ clknet_leaf_29_clk _0713_ VGND VGND VPWR VPWR rf.registers\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6765_ _3296_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7148__S _3455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8504_ net453 net33 _4227_ VGND VGND VPWR VPWR _4235_ sky130_fd_sc_hd__mux2_1
X_5716_ _2387_ _2393_ _1146_ VGND VGND VPWR VPWR _2469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9484_ clknet_leaf_50_clk _0644_ VGND VGND VPWR VPWR rf.registers\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6696_ net485 _3002_ _3253_ VGND VGND VPWR VPWR _3260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8435_ _4198_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _1168_ _1821_ _2401_ VGND VGND VPWR VPWR _2402_ sky130_fd_sc_hd__o21ba_1
XANTENNA__7672__A _3771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8366_ net475 _3442_ _4155_ VGND VGND VPWR VPWR _4162_ sky130_fd_sc_hd__mux2_1
X_5578_ _2331_ _2332_ _2333_ VGND VGND VPWR VPWR _2334_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4440__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold230 rf.registers\[14\]\[12\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold241 rf.registers\[7\]\[8\] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
X_7317_ _3050_ net733 _3602_ VGND VGND VPWR VPWR _3606_ sky130_fd_sc_hd__mux2_1
Xhold252 rf.registers\[5\]\[5\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _1283_ _1284_ _1198_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__mux2_1
X_8297_ _4125_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__clkbuf_1
Xhold263 rf.registers\[2\]\[14\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 rf.registers\[8\]\[7\] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4300__S _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold285 rf.registers\[25\]\[14\] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 rf.registers\[6\]\[2\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7248_ _3569_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
X_7179_ net637 _3483_ _3528_ VGND VGND VPWR VPWR _3532_ sky130_fd_sc_hd__mux2_1
XANTENNA__7611__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6751__A _3266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8442__S _4168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4271__A _1026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5208__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6897__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 A3[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4446__A _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4880_ _1512_ net96 _1635_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__and3_1
XANTENNA__5447__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6550_ net683 _3139_ _3179_ VGND VGND VPWR VPWR _3182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5501_ rf.registers\[16\]\[6\] rf.registers\[17\]\[6\] rf.registers\[18\]\[6\] rf.registers\[19\]\[6\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4670__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6481_ net30 VGND VGND VPWR VPWR _3143_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_125_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8220_ net948 _3500_ _4083_ VGND VGND VPWR VPWR _4085_ sky130_fd_sc_hd__mux2_1
X_5432_ _1686_ _2185_ _2187_ _1699_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5363_ rf.registers\[4\]\[15\] rf.registers\[5\]\[15\] rf.registers\[6\]\[15\] rf.registers\[7\]\[15\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__mux4_1
X_8151_ _4048_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5216__S _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7102_ net335 _3485_ _3477_ VGND VGND VPWR VPWR _3486_ sky130_fd_sc_hd__mux2_1
X_4314_ _1064_ _1069_ _1037_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5294_ _1673_ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__buf_4
X_8082_ net891 _3497_ _4011_ VGND VGND VPWR VPWR _4012_ sky130_fd_sc_hd__mux2_1
X_7033_ _3439_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8527__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7431__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8984_ clknet_leaf_11_clk _0144_ VGND VGND VPWR VPWR rf.registers\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6252__A1 _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7935_ _3933_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8262__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7866_ _3124_ net655 _3891_ VGND VGND VPWR VPWR _3897_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_60_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6817_ _3324_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7797_ _3860_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9536_ clknet_leaf_70_clk _0696_ VGND VGND VPWR VPWR rf.registers\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5763__B1 _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6748_ _3287_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4661__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9467_ clknet_leaf_26_clk _0627_ VGND VGND VPWR VPWR rf.registers\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6679_ net560 _3130_ _3242_ VGND VGND VPWR VPWR _3251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5915__A _1464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6510__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8418_ _4189_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9398_ clknet_leaf_33_clk _0558_ VGND VGND VPWR VPWR rf.registers\[24\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8349_ net494 _3493_ _4144_ VGND VGND VPWR VPWR _4153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6491__A1 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6481__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8172__S _4024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_28_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5429__S0 _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5097__A _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4652__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7516__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6420__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7259__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8347__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7251__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6234__A1 _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5981_ _2571_ _2605_ _2720_ _1087_ _2721_ VGND VGND VPWR VPWR _2722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7720_ _3043_ net518 _3819_ VGND VGND VPWR VPWR _3820_ sky130_fd_sc_hd__mux2_1
XANTENNA__8082__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4340__S0 _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4932_ rf.registers\[28\]\[23\] rf.registers\[29\]\[23\] rf.registers\[30\]\[23\]
+ rf.registers\[31\]\[23\] _1676_ _1681_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_44_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7651_ _3771_ VGND VGND VPWR VPWR _3783_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__5719__B _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4863_ rf.registers\[20\]\[18\] rf.registers\[21\]\[18\] rf.registers\[22\]\[18\]
+ rf.registers\[23\]\[18\] net109 _1202_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6602_ _3210_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_103_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_14 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7582_ _3746_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
X_4794_ rf.registers\[8\]\[10\] rf.registers\[9\]\[10\] rf.registers\[10\]\[10\] rf.registers\[11\]\[10\]
+ net117 _1053_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__mux4_1
X_9321_ clknet_leaf_51_clk _0481_ VGND VGND VPWR VPWR rf.registers\[21\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6533_ net443 _3122_ _3168_ VGND VGND VPWR VPWR _3173_ sky130_fd_sc_hd__mux2_1
XANTENNA__5735__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6330__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9252_ clknet_leaf_48_clk _0412_ VGND VGND VPWR VPWR rf.registers\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6464_ _3131_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8203_ net154 _3483_ _4072_ VGND VGND VPWR VPWR _4076_ sky130_fd_sc_hd__mux2_1
X_5415_ rf.registers\[4\]\[12\] rf.registers\[5\]\[12\] rf.registers\[6\]\[12\] rf.registers\[7\]\[12\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2171_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9183_ clknet_leaf_74_clk _0343_ VGND VGND VPWR VPWR rf.registers\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6395_ _3083_ net1126 _3065_ VGND VGND VPWR VPWR _3084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8134_ _4039_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__clkbuf_1
X_5346_ _1060_ _2101_ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__nand2_4
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8065_ net519 _3481_ _4000_ VGND VGND VPWR VPWR _4003_ sky130_fd_sc_hd__mux2_1
X_5277_ _1777_ _2024_ _2032_ VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__a21oi_4
XANTENNA__6473__A1 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7016_ _3430_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5681__C1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8967_ clknet_leaf_66_clk _0127_ VGND VGND VPWR VPWR rf.registers\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7918_ _3924_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__clkbuf_1
X_8898_ clknet_leaf_54_clk _0058_ VGND VGND VPWR VPWR rf.registers\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7849_ _3107_ net604 _3880_ VGND VGND VPWR VPWR _3888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4634__S1 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9519_ clknet_leaf_8_clk _0679_ VGND VGND VPWR VPWR rf.registers\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7336__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8150__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4398__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4695__S _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7071__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4570__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4625__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput12 A3[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
Xinput23 WD3[18] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput34 WD3[28] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput45 WD3[9] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold807 rf.registers\[25\]\[10\] VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8141__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold818 rf.registers\[11\]\[4\] VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 rf.registers\[7\]\[21\] VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5050__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5200_ _1954_ _1955_ _1889_ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6180_ _2866_ _2909_ _2327_ VGND VGND VPWR VPWR _2910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5711__A_N _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5131_ rf.registers\[16\]\[31\] rf.registers\[17\]\[31\] rf.registers\[18\]\[31\]
+ rf.registers\[19\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__mux4_1
XANTENNA__8077__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5062_ _1816_ _1817_ _1686_ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_6__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8821_ clknet_leaf_32_clk _1005_ VGND VGND VPWR VPWR rf.registers\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7955__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8752_ clknet_leaf_13_clk _0936_ VGND VGND VPWR VPWR rf.registers\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_5964_ _2549_ _2705_ _2104_ VGND VGND VPWR VPWR _2706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7703_ _3027_ net1019 _3808_ VGND VGND VPWR VPWR _3811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4915_ _1670_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__clkbuf_8
X_8683_ clknet_leaf_4_clk _0867_ VGND VGND VPWR VPWR rf.registers\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5895_ _1572_ _2595_ _2639_ VGND VGND VPWR VPWR _2640_ sky130_fd_sc_hd__nand3_1
XFILLER_0_114_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5718__A0 _2469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7634_ _3774_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4846_ _1587_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7565_ _3025_ net690 _3736_ VGND VGND VPWR VPWR _3738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4777_ _1529_ _1530_ _1531_ _1532_ _1040_ _1038_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__mux4_2
XFILLER_0_105_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7156__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9304_ clknet_leaf_27_clk _0464_ VGND VGND VPWR VPWR rf.registers\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6516_ net231 _3105_ _3157_ VGND VGND VPWR VPWR _3164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7496_ _3701_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_151_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9235_ clknet_leaf_34_clk _0395_ VGND VGND VPWR VPWR rf.registers\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6447_ net18 VGND VGND VPWR VPWR _3120_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6694__A1 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9166_ clknet_leaf_29_clk _0326_ VGND VGND VPWR VPWR rf.registers\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6378_ _3072_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__clkbuf_1
X_8117_ _4030_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__clkbuf_1
X_5329_ rf.registers\[28\]\[1\] rf.registers\[29\]\[1\] rf.registers\[30\]\[1\] rf.registers\[31\]\[1\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__mux4_1
X_9097_ clknet_leaf_50_clk _0257_ VGND VGND VPWR VPWR rf.registers\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8048_ net649 _3464_ _3989_ VGND VGND VPWR VPWR _3994_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__S0 _1267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8199__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5118__A1_N _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7855__A _3879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8450__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5185__B2 _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4719__A _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4791__S0 _1041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5314__S _1645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4327__A1_N _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5099__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4700_ rf.registers\[4\]\[12\] rf.registers\[5\]\[12\] rf.registers\[6\]\[12\] rf.registers\[7\]\[12\]
+ net1161 _1279_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8360__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5680_ _1148_ _2432_ _2433_ _2337_ VGND VGND VPWR VPWR _2434_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4631_ rf.registers\[28\]\[6\] rf.registers\[29\]\[6\] rf.registers\[30\]\[6\] rf.registers\[31\]\[6\]
+ net100 _1221_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5271__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7350_ _3083_ net1000 _3613_ VGND VGND VPWR VPWR _3623_ sky130_fd_sc_hd__mux2_1
X_4562_ rf.registers\[16\]\[31\] rf.registers\[17\]\[31\] rf.registers\[18\]\[31\]
+ rf.registers\[19\]\[31\] _1200_ _1202_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6301_ net14 VGND VGND VPWR VPWR _3019_ sky130_fd_sc_hd__clkbuf_2
Xhold604 rf.registers\[10\]\[1\] VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold615 rf.registers\[8\]\[9\] VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 rf.registers\[5\]\[4\] VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__dlygate4sd3_1
X_7281_ _3586_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_133_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4493_ rf.registers\[12\]\[20\] rf.registers\[13\]\[20\] rf.registers\[14\]\[20\]
+ rf.registers\[15\]\[20\] _1201_ _1203_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__mux4_1
Xhold637 rf.registers\[22\]\[19\] VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 rf.registers\[29\]\[12\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__dlygate4sd3_1
X_9020_ clknet_leaf_12_clk _0180_ VGND VGND VPWR VPWR rf.registers\[31\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold659 rf.registers\[21\]\[4\] VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _2923_ _2384_ _1148_ VGND VGND VPWR VPWR _2959_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6163_ _2887_ _2893_ VGND VGND VPWR VPWR _2894_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4782__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4629__A _1370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5114_ rf.registers\[4\]\[16\] rf.registers\[5\]\[16\] rf.registers\[6\]\[16\] rf.registers\[7\]\[16\]
+ _1822_ _1823_ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__mux4_1
X_6094_ net134 _2828_ VGND VGND VPWR VPWR _2829_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8535__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5045_ _1758_ _1798_ _1800_ VGND VGND VPWR VPWR _1801_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8804_ clknet_leaf_51_clk _0988_ VGND VGND VPWR VPWR rf.registers\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6055__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6996_ net203 _3105_ _3413_ VGND VGND VPWR VPWR _3420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4837__S1 _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8735_ clknet_leaf_73_clk _0919_ VGND VGND VPWR VPWR rf.registers\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5947_ _2689_ _2669_ net1166 VGND VGND VPWR VPWR _2690_ sky130_fd_sc_hd__and3b_1
XFILLER_0_149_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8666_ clknet_leaf_21_clk _0850_ VGND VGND VPWR VPWR rf.registers\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5878_ _2623_ VGND VGND VPWR VPWR _2624_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone26 A2[0] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_16
XANTENNA__6364__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7617_ _3077_ net568 _3758_ VGND VGND VPWR VPWR _3765_ sky130_fd_sc_hd__mux2_1
X_4829_ _1583_ _1584_ _1036_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8597_ clknet_leaf_31_clk _0781_ VGND VGND VPWR VPWR rf.registers\[22\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5195__A _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5262__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7548_ _3728_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6116__B1 _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7479_ _3075_ net1072 _3686_ VGND VGND VPWR VPWR _3692_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7864__A0 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5014__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9218_ clknet_leaf_60_clk _0378_ VGND VGND VPWR VPWR rf.registers\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9149_ clknet_leaf_3_clk _0309_ VGND VGND VPWR VPWR rf.registers\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4773__S0 _1290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4525__S0 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4828__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8180__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6355__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7524__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output78_A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4764__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__A _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5979__S _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6850_ _3342_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5801_ _2254_ _2425_ _2431_ _2337_ VGND VGND VPWR VPWR _2551_ sky130_fd_sc_hd__o22a_1
XANTENNA__4819__S1 _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6781_ net235 _3095_ _3304_ VGND VGND VPWR VPWR _3306_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8090__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8520_ rf.registers\[10\]\[3\] net39 _3007_ VGND VGND VPWR VPWR _4243_ sky130_fd_sc_hd__mux2_1
X_5732_ _2482_ _2484_ VGND VGND VPWR VPWR _2485_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6603__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4912__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8335__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8451_ _4207_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5663_ _1662_ VGND VGND VPWR VPWR _2417_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7402_ _3651_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5244__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4614_ _1171_ _1359_ _1365_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_154_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8382_ net557 _3458_ _4169_ VGND VGND VPWR VPWR _4171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5594_ _1758_ _2175_ _1839_ VGND VGND VPWR VPWR _2349_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7333_ _3614_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
Xhold401 rf.registers\[22\]\[20\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4545_ rf.registers\[16\]\[27\] rf.registers\[17\]\[27\] rf.registers\[18\]\[27\]
+ rf.registers\[19\]\[27\] _1262_ _1263_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__mux4_2
XFILLER_0_4_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold412 rf.registers\[16\]\[18\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold423 rf.registers\[27\]\[7\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5743__A _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold434 rf.registers\[5\]\[23\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 rf.registers\[13\]\[11\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7264_ _3064_ net635 _3577_ VGND VGND VPWR VPWR _3578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold456 rf.registers\[30\]\[23\] VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _1199_ _1231_ _1213_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__a21o_1
Xhold467 rf.registers\[4\]\[0\] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
X_9003_ clknet_leaf_2_clk _0163_ VGND VGND VPWR VPWR rf.registers\[31\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold478 rf.registers\[8\]\[18\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 rf.registers\[2\]\[29\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _1962_ _2942_ _2421_ VGND VGND VPWR VPWR _2943_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7195_ _3540_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _2808_ _2830_ _2840_ _2854_ VGND VGND VPWR VPWR _2878_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_51_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7074__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8271__A0 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4793__S _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8265__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6077_ _2601_ VGND VGND VPWR VPWR _2813_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_146_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6821__A1 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5028_ rf.registers\[16\]\[20\] rf.registers\[17\]\[20\] rf.registers\[18\]\[20\]
+ rf.registers\[19\]\[20\] _1782_ _1680_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__mux4_1
XANTENNA__5180__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8023__A0 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6979_ net1023 _3017_ _3375_ VGND VGND VPWR VPWR _3410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5918__A _2175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7609__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5483__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8718_ clknet_leaf_29_clk _0902_ VGND VGND VPWR VPWR rf.registers\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8326__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6337__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8649_ clknet_leaf_47_clk _0833_ VGND VGND VPWR VPWR rf.registers\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5235__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4994__S0 _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7344__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7837__A0 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5653__A _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold990 rf.registers\[25\]\[25\] VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5799__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8262__A0 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6484__A net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6812__A1 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5171__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6423__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5226__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4985__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4330_ _1060_ _1085_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6000_ _2584_ _2731_ _2736_ _2496_ _2739_ VGND VGND VPWR VPWR _2740_ sky130_fd_sc_hd__a221o_1
XANTENNA__6394__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4907__A _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5502__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7951_ net1082 _3504_ _3938_ VGND VGND VPWR VPWR _3942_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6902_ _3369_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__clkbuf_1
X_7882_ _3905_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8556__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6833_ net424 _3002_ _3326_ VGND VGND VPWR VPWR _3333_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7429__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6333__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5465__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9552_ clknet_leaf_13_clk _0712_ VGND VGND VPWR VPWR rf.registers\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6764_ _3077_ net593 _3289_ VGND VGND VPWR VPWR _3296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8503_ _4234_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__clkbuf_1
X_5715_ _1666_ VGND VGND VPWR VPWR _2468_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9483_ clknet_leaf_5_clk _0643_ VGND VGND VPWR VPWR rf.registers\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6695_ _3259_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8434_ net1036 net32 _4191_ VGND VGND VPWR VPWR _4198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5646_ net82 _1859_ VGND VGND VPWR VPWR _2401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8365_ _4161_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__clkbuf_1
X_5577_ net48 VGND VGND VPWR VPWR _2333_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__7164__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold220 rf.registers\[13\]\[31\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7316_ _3605_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
Xhold231 rf.registers\[20\]\[1\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ rf.registers\[24\]\[26\] rf.registers\[25\]\[26\] rf.registers\[26\]\[26\]
+ rf.registers\[27\]\[26\] net1155 _1183_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__mux4_2
Xhold242 rf.registers\[24\]\[14\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
X_8296_ _3145_ net404 _4119_ VGND VGND VPWR VPWR _4125_ sky130_fd_sc_hd__mux2_1
Xhold253 rf.registers\[3\]\[14\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 rf.registers\[7\]\[0\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold275 rf.registers\[25\]\[0\] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4728__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7247_ _3048_ net730 _3566_ VGND VGND VPWR VPWR _3569_ sky130_fd_sc_hd__mux2_1
Xhold286 rf.registers\[13\]\[10\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _1025_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__clkbuf_8
Xhold297 rf.registers\[5\]\[19\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
X_7178_ _3531_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
X_6129_ _2496_ _2859_ _2861_ _2504_ VGND VGND VPWR VPWR _2862_ sky130_fd_sc_hd__a211o_1
XANTENNA__6508__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5153__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4900__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6243__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clone22_A _1172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5781__A1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5781__B2 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5208__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4698__S _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5533__A1 _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7074__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7802__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5392__S0 _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5322__S _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5144__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7249__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7210__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5447__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5221__B1 _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5500_ rf.registers\[20\]\[6\] rf.registers\[21\]\[6\] rf.registers\[22\]\[6\] rf.registers\[23\]\[6\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6480_ _3142_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5431_ _1711_ _2186_ VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8150_ net817 _3497_ _4047_ VGND VGND VPWR VPWR _4048_ sky130_fd_sc_hd__mux2_1
X_5362_ _1678_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7101_ net19 VGND VGND VPWR VPWR _3485_ sky130_fd_sc_hd__buf_2
X_4313_ _1067_ _1068_ _1035_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8081_ _3988_ VGND VGND VPWR VPWR _4011_ sky130_fd_sc_hd__clkbuf_8
X_5293_ _2045_ _2048_ _1696_ VGND VGND VPWR VPWR _2049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7032_ net498 _3141_ _3435_ VGND VGND VPWR VPWR _3439_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5135__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8983_ clknet_leaf_34_clk _0143_ VGND VGND VPWR VPWR rf.registers\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_7934_ net664 _3487_ _3927_ VGND VGND VPWR VPWR _3933_ sky130_fd_sc_hd__mux2_1
XANTENNA__8529__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7865_ _3896_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5468__A _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4372__A _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6816_ net444 _3130_ _3315_ VGND VGND VPWR VPWR _3324_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7796_ net395 _3485_ _3855_ VGND VGND VPWR VPWR _3860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5187__B _1942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9535_ clknet_leaf_71_clk _0695_ VGND VGND VPWR VPWR rf.registers\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6998__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5763__A1 _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6747_ _3060_ net575 _3278_ VGND VGND VPWR VPWR _3287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9466_ clknet_leaf_18_clk _0626_ VGND VGND VPWR VPWR rf.registers\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6678_ _3250_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5915__B _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8417_ net529 _3493_ _4180_ VGND VGND VPWR VPWR _4189_ sky130_fd_sc_hd__mux2_1
X_5629_ _1799_ _1979_ VGND VGND VPWR VPWR _2384_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_154_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9397_ clknet_leaf_31_clk _0557_ VGND VGND VPWR VPWR rf.registers\[24\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8348_ _4152_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8279_ _3128_ net446 _4108_ VGND VGND VPWR VPWR _4116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5429__S1 _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4282__A _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7532__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output60_A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4457__A _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6219__C1 _1085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5980_ _2468_ _2530_ _2426_ _2472_ _2503_ VGND VGND VPWR VPWR _2721_ sky130_fd_sc_hd__a41o_1
XFILLER_0_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4931_ _1682_ _1683_ _1686_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__mux2_1
XANTENNA__5993__A1 _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4340__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5288__A _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7650_ _3782_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4862_ _1239_ _1609_ _1617_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6601_ _3050_ net572 _3206_ VGND VGND VPWR VPWR _3210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_15 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7581_ _3041_ net1030 _3736_ VGND VGND VPWR VPWR _3746_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4793_ _1545_ _1548_ _1037_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7707__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9320_ clknet_leaf_48_clk _0480_ VGND VGND VPWR VPWR rf.registers\[21\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6611__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ _3172_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4920__A _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9251_ clknet_leaf_68_clk _0411_ VGND VGND VPWR VPWR rf.registers\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5735__B _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6463_ net280 _3130_ _3114_ VGND VGND VPWR VPWR _3131_ sky130_fd_sc_hd__mux2_1
XANTENNA__5227__S _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8202_ _4075_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5414_ _1699_ _2169_ VGND VGND VPWR VPWR _2170_ sky130_fd_sc_hd__nand2_1
X_9182_ clknet_leaf_74_clk _0342_ VGND VGND VPWR VPWR rf.registers\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6170__A1 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6394_ net35 VGND VGND VPWR VPWR _3083_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8133_ net624 _3481_ _4036_ VGND VGND VPWR VPWR _4039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5345_ _1664_ _1084_ VGND VGND VPWR VPWR _2101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5751__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8064_ _4002_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__clkbuf_1
X_5276_ _2026_ _2028_ _2031_ _1766_ _1672_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__o221a_1
X_7015_ net654 _3124_ _3424_ VGND VGND VPWR VPWR _3430_ sky130_fd_sc_hd__mux2_1
XANTENNA__7670__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5108__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8273__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8966_ clknet_leaf_0_clk _0126_ VGND VGND VPWR VPWR rf.registers\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7917_ net416 _3470_ _3916_ VGND VGND VPWR VPWR _3924_ sky130_fd_sc_hd__mux2_1
X_8897_ clknet_leaf_57_clk _0057_ VGND VGND VPWR VPWR rf.registers\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7848_ _3887_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5736__A1 _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7779_ net369 _3468_ _3844_ VGND VGND VPWR VPWR _3851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7617__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9518_ clknet_leaf_29_clk _0678_ VGND VGND VPWR VPWR rf.registers\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9449_ clknet_leaf_65_clk _0609_ VGND VGND VPWR VPWR rf.registers\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5137__S _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4398__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8448__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7352__S _3590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4570__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 A3[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput24 WD3[19] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput35 WD3[29] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput46 WE3 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_4
XFILLER_0_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold808 rf.registers\[28\]\[10\] VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold819 rf.registers\[13\]\[24\] VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8358__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5130_ rf.registers\[28\]\[31\] rf.registers\[29\]\[31\] rf.registers\[30\]\[31\]
+ rf.registers\[31\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5338__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7652__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5061_ rf.registers\[0\]\[18\] rf.registers\[1\]\[18\] rf.registers\[2\]\[18\] rf.registers\[3\]\[18\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8820_ clknet_leaf_30_clk _1004_ VGND VGND VPWR VPWR rf.registers\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4915__A _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5963_ _2624_ _2704_ _2501_ VGND VGND VPWR VPWR _2705_ sky130_fd_sc_hd__mux2_1
X_8751_ clknet_leaf_11_clk _0935_ VGND VGND VPWR VPWR rf.registers\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7702_ _3810_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4914_ _1640_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__clkbuf_4
X_5894_ _2638_ net121 _2593_ _2594_ VGND VGND VPWR VPWR _2639_ sky130_fd_sc_hd__or4_4
X_8682_ clknet_leaf_7_clk _0866_ VGND VGND VPWR VPWR rf.registers\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7633_ net652 _3458_ _3772_ VGND VGND VPWR VPWR _3774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5718__A1 _2470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4845_ _1215_ _1592_ _1596_ _1600_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_28_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7437__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7564_ _3737_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
X_4776_ rf.registers\[24\]\[9\] rf.registers\[25\]\[9\] rf.registers\[26\]\[9\] rf.registers\[27\]\[9\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__mux4_2
XFILLER_0_117_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6515_ _3163_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9303_ clknet_leaf_33_clk _0463_ VGND VGND VPWR VPWR rf.registers\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7495_ _3019_ net551 _3700_ VGND VGND VPWR VPWR _3701_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7340__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6446_ _3119_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__clkbuf_1
X_9234_ clknet_leaf_27_clk _0394_ VGND VGND VPWR VPWR rf.registers\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4796__S _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9165_ clknet_leaf_44_clk _0325_ VGND VGND VPWR VPWR rf.registers\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6377_ _3071_ net1012 _3065_ VGND VGND VPWR VPWR _3072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_27_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8116_ net542 _3464_ _4025_ VGND VGND VPWR VPWR _4030_ sky130_fd_sc_hd__mux2_1
X_5328_ rf.registers\[24\]\[1\] rf.registers\[25\]\[1\] rf.registers\[26\]\[1\] rf.registers\[27\]\[1\]
+ _1673_ _1690_ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__mux4_1
XANTENNA__5329__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9096_ clknet_leaf_49_clk _0256_ VGND VGND VPWR VPWR rf.registers\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8047_ _3993_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7643__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5259_ _1777_ _2006_ _2010_ _2014_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_54_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6516__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5501__S0 _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8949_ clknet_leaf_25_clk _0109_ VGND VGND VPWR VPWR rf.registers\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_rebuffer32_A _1528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6134__A1 _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8178__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4791__S1 _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6426__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7398__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload5_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7257__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4630_ rf.registers\[24\]\[6\] rf.registers\[25\]\[6\] rf.registers\[26\]\[6\] rf.registers\[27\]\[6\]
+ _1219_ _1221_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__mux4_2
XFILLER_0_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4561_ rf.registers\[20\]\[31\] rf.registers\[21\]\[31\] rf.registers\[22\]\[31\]
+ rf.registers\[23\]\[31\] net109 _1202_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6300_ _3018_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold605 rf.registers\[16\]\[8\] VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7280_ _3081_ net678 _3577_ VGND VGND VPWR VPWR _3586_ sky130_fd_sc_hd__mux2_1
XANTENNA__5559__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold616 rf.registers\[1\]\[8\] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4492_ _1190_ _1247_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_133_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold627 rf.registers\[0\]\[20\] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 rf.registers\[23\]\[10\] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6231_ _2380_ _2383_ VGND VGND VPWR VPWR _2958_ sky130_fd_sc_hd__or2b_1
Xhold649 rf.registers\[23\]\[26\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8088__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6397__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5505__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6162_ _2891_ _2892_ VGND VGND VPWR VPWR _2893_ sky130_fd_sc_hd__or2_1
XANTENNA__4782__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4629__B _1384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5113_ _1717_ _1868_ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__nor2_1
X_6093_ _1512_ net105 net1160 _2658_ _2741_ VGND VGND VPWR VPWR _2828_ sky130_fd_sc_hd__a41o_1
XANTENNA__7720__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5044_ _1799_ VGND VGND VPWR VPWR _1800_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8803_ clknet_leaf_54_clk _0987_ VGND VGND VPWR VPWR rf.registers\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8050__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5939__A1 _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6995_ _3419_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4298__S0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8734_ clknet_leaf_72_clk _0918_ VGND VGND VPWR VPWR rf.registers\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_5946_ _2687_ _2688_ VGND VGND VPWR VPWR _2689_ sky130_fd_sc_hd__or2_4
XFILLER_0_125_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5877_ _2581_ _2622_ _1146_ VGND VGND VPWR VPWR _2623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8665_ clknet_leaf_20_clk _0849_ VGND VGND VPWR VPWR rf.registers\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4828_ rf.registers\[0\]\[16\] rf.registers\[1\]\[16\] rf.registers\[2\]\[16\] rf.registers\[3\]\[16\]
+ net1158 _1183_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__mux4_1
X_7616_ _3764_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
Xclone27 _1027_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone38 _1065_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_16
X_8596_ clknet_leaf_42_clk _0780_ VGND VGND VPWR VPWR rf.registers\[22\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4759_ _1513_ _1514_ _1035_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__mux2_1
X_7547_ _3075_ net721 _3722_ VGND VGND VPWR VPWR _3728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4470__S0 _1220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7313__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7478_ _3691_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
X_9217_ clknet_leaf_60_clk _0377_ VGND VGND VPWR VPWR rf.registers\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_56_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6429_ net627 _3107_ _3093_ VGND VGND VPWR VPWR _3108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9148_ clknet_leaf_12_clk _0308_ VGND VGND VPWR VPWR rf.registers\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4773__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9079_ clknet_leaf_34_clk _0239_ VGND VGND VPWR VPWR rf.registers\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4525__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6246__S _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4289__S0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7077__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5386__A _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4290__A _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4764__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4465__A _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5800_ _2439_ _2424_ _2501_ VGND VGND VPWR VPWR _2550_ sky130_fd_sc_hd__mux2_1
X_6780_ _3305_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5731_ _2449_ _2451_ _2483_ VGND VGND VPWR VPWR _2484_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5296__A _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4404__S _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8450_ net623 net25 _4205_ VGND VGND VPWR VPWR _4207_ sky130_fd_sc_hd__mux2_1
X_5662_ _2376_ _2407_ _2408_ _2416_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_154_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7401_ _3064_ net971 _3650_ VGND VGND VPWR VPWR _3651_ sky130_fd_sc_hd__mux2_1
X_4613_ _1214_ _1368_ _1239_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__o21ai_1
X_8381_ _4170_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__clkbuf_1
X_5593_ _2343_ _2346_ _2347_ VGND VGND VPWR VPWR _2348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5102__A1_N _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7715__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7332_ _3064_ net1079 _3613_ VGND VGND VPWR VPWR _3614_ sky130_fd_sc_hd__mux2_1
X_4544_ rf.registers\[20\]\[27\] rf.registers\[21\]\[27\] rf.registers\[22\]\[27\]
+ rf.registers\[23\]\[27\] _1262_ _1263_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold402 rf.registers\[3\]\[25\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8400__A _4168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold413 rf.registers\[15\]\[2\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold424 rf.registers\[3\]\[0\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
X_7263_ _3554_ VGND VGND VPWR VPWR _3577_ sky130_fd_sc_hd__clkbuf_8
Xhold435 rf.registers\[31\]\[27\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 rf.registers\[3\]\[4\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ rf.registers\[0\]\[28\] rf.registers\[1\]\[28\] rf.registers\[2\]\[28\] rf.registers\[3\]\[28\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__mux4_1
Xhold457 rf.registers\[7\]\[20\] VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 rf.registers\[25\]\[5\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9002_ clknet_leaf_45_clk _0162_ VGND VGND VPWR VPWR rf.registers\[31\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6214_ _2426_ _2591_ VGND VGND VPWR VPWR _2942_ sky130_fd_sc_hd__nand2_1
Xhold479 rf.registers\[3\]\[1\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7194_ net539 _3497_ _3539_ VGND VGND VPWR VPWR _3540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _2875_ _2876_ VGND VGND VPWR VPWR _2877_ sky130_fd_sc_hd__or2_1
XANTENNA__8546__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7450__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _2773_ _2809_ _2810_ _2811_ VGND VGND VPWR VPWR _2812_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_146_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5085__A1 _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ rf.registers\[20\]\[20\] rf.registers\[21\]\[20\] rf.registers\[22\]\[20\]
+ rf.registers\[23\]\[20\] _1782_ _1680_ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__mux4_1
XANTENNA__5180__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4388__A1_N _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8281__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6978_ _3409_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8717_ clknet_leaf_44_clk _0901_ VGND VGND VPWR VPWR rf.registers\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5929_ _2547_ _2672_ _1147_ VGND VGND VPWR VPWR _2673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4314__S _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8648_ clknet_leaf_63_clk _0832_ VGND VGND VPWR VPWR rf.registers\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7534__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8579_ clknet_leaf_68_clk _0763_ VGND VGND VPWR VPWR rf.registers\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7625__S _3735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4994__S1 _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5848__B1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold980 rf.registers\[27\]\[27\] VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 rf.registers\[26\]\[2\] VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4520__B1 _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4984__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8456__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5171__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6704__S _3230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4587__B1 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4682__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4985__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5055__S _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4894__S net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8366__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7270__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7950_ _3941_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6901_ net545 _3002_ _3362_ VGND VGND VPWR VPWR _3369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7881_ _3139_ net713 _3902_ VGND VGND VPWR VPWR _3905_ sky130_fd_sc_hd__mux2_1
XANTENNA__4923__A _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6832_ _3332_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9551_ clknet_leaf_11_clk _0711_ VGND VGND VPWR VPWR rf.registers\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6763_ _3295_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8502_ net660 net32 _4227_ VGND VGND VPWR VPWR _4234_ sky130_fd_sc_hd__mux2_1
XANTENNA__7516__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5714_ _2105_ _2462_ _2466_ VGND VGND VPWR VPWR _2467_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9482_ clknet_leaf_63_clk _0642_ VGND VGND VPWR VPWR rf.registers\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6694_ net612 _3145_ _3253_ VGND VGND VPWR VPWR _3259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8433_ _4197_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5645_ _2398_ _2399_ VGND VGND VPWR VPWR _2400_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7445__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5754__A _1125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5576_ _1669_ _1660_ VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8364_ net956 _3508_ _4155_ VGND VGND VPWR VPWR _4161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold210 rf.registers\[6\]\[28\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7819__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold221 rf.registers\[3\]\[3\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
X_7315_ _3048_ net534 _3602_ VGND VGND VPWR VPWR _3605_ sky130_fd_sc_hd__mux2_1
X_4527_ rf.registers\[28\]\[26\] rf.registers\[29\]\[26\] rf.registers\[30\]\[26\]
+ rf.registers\[31\]\[26\] net1155 _1183_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold232 rf.registers\[17\]\[6\] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
X_8295_ _4124_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__clkbuf_1
Xhold243 rf.registers\[18\]\[28\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold254 rf.registers\[12\]\[30\] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8492__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold265 rf.registers\[10\]\[10\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7246_ _3568_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
Xhold276 rf.registers\[9\]\[26\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ _1213_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold287 rf.registers\[9\]\[6\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4728__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold298 rf.registers\[24\]\[30\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
X_7177_ net232 _3481_ _3528_ VGND VGND VPWR VPWR _3531_ sky130_fd_sc_hd__mux2_1
X_4389_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__clkbuf_4
X_6128_ _2373_ _2572_ _2823_ _2569_ _2860_ VGND VGND VPWR VPWR _2861_ sky130_fd_sc_hd__a221o_1
XANTENNA__4817__B _1542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _2102_ _2488_ VGND VGND VPWR VPWR _2795_ sky130_fd_sc_hd__nor2_1
XANTENNA__5153__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4900__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4664__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8483__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8186__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5392__S1 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7090__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6797__A1 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7994__A0 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5144__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5221__A1 _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4655__S0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4407__S0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5430_ rf.registers\[8\]\[11\] rf.registers\[9\]\[11\] rf.registers\[10\]\[11\] rf.registers\[11\]\[11\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6182__C1 _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5361_ _1702_ VGND VGND VPWR VPWR _2117_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4312_ rf.registers\[24\]\[5\] rf.registers\[25\]\[5\] rf.registers\[26\]\[5\] rf.registers\[27\]\[5\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7100_ _3484_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8080_ _4010_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__clkbuf_1
X_5292_ _2046_ _2047_ _2044_ VGND VGND VPWR VPWR _2048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7031_ _3438_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8096__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4918__A _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6609__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5513__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8982_ clknet_leaf_33_clk _0142_ VGND VGND VPWR VPWR rf.registers\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7985__A0 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5135__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7933_ _3932_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5749__A _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7864_ _3122_ net739 _3891_ VGND VGND VPWR VPWR _3896_ sky130_fd_sc_hd__mux2_1
XANTENNA__6571__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6815_ _3323_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4372__B _1127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7795_ _3859_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9534_ clknet_leaf_72_clk _0694_ VGND VGND VPWR VPWR rf.registers\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6746_ _3286_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9465_ clknet_leaf_19_clk _0625_ VGND VGND VPWR VPWR rf.registers\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6677_ net643 _3128_ _3242_ VGND VGND VPWR VPWR _3250_ sky130_fd_sc_hd__mux2_1
XANTENNA__7175__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8416_ _4188_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5628_ _1668_ _1959_ VGND VGND VPWR VPWR _2383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9396_ clknet_leaf_42_clk _0556_ VGND VGND VPWR VPWR rf.registers\[24\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_154_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5071__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4723__B1 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8347_ net622 _3491_ _4144_ VGND VGND VPWR VPWR _4152_ sky130_fd_sc_hd__mux2_1
X_5559_ rf.registers\[8\]\[5\] rf.registers\[9\]\[5\] rf.registers\[10\]\[5\] rf.registers\[11\]\[5\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__mux4_1
XANTENNA__7903__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8278_ _4115_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__clkbuf_1
X_7229_ _3559_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5423__S _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5659__A _2097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7728__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4637__S0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7813__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8456__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6429__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output53_A net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5569__A _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4930_ _1685_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__buf_4
X_4861_ _1611_ _1613_ _1616_ _1214_ _1170_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__a221o_1
X_6600_ _3209_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7580_ _3745_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4792_ _1546_ _1547_ _1034_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__mux2_1
XANTENNA_16 _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6942__A1 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6531_ net149 _3120_ _3168_ VGND VGND VPWR VPWR _3172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9250_ clknet_leaf_58_clk _0410_ VGND VGND VPWR VPWR rf.registers\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6462_ net23 VGND VGND VPWR VPWR _3130_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5053__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8201_ net363 _3481_ _4072_ VGND VGND VPWR VPWR _4075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5413_ _2167_ _2168_ _1711_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9181_ clknet_leaf_15_clk _0341_ VGND VGND VPWR VPWR rf.registers\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6393_ _3082_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__clkbuf_1
X_5344_ _2083_ _2099_ _1148_ VGND VGND VPWR VPWR _2100_ sky130_fd_sc_hd__mux2_1
X_8132_ _4038_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8063_ net898 _3479_ _4000_ VGND VGND VPWR VPWR _4002_ sky130_fd_sc_hd__mux2_1
X_5275_ _2029_ _2030_ _1901_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7014_ _3429_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5681__A1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8554__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5108__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8965_ clknet_leaf_62_clk _0125_ VGND VGND VPWR VPWR rf.registers\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4383__A _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7916_ _3923_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__clkbuf_1
X_8896_ clknet_leaf_60_clk _0056_ VGND VGND VPWR VPWR rf.registers\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7847_ _3105_ net481 _3880_ VGND VGND VPWR VPWR _3887_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4619__S0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5197__B1 _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6802__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7778_ _3850_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6933__A1 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9517_ clknet_leaf_29_clk _0677_ VGND VGND VPWR VPWR rf.registers\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6729_ _3277_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9448_ clknet_leaf_63_clk _0608_ VGND VGND VPWR VPWR rf.registers\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9379_ clknet_leaf_67_clk _0539_ VGND VGND VPWR VPWR rf.registers\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7633__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5942__A _1464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8464__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4858__S0 _1173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6712__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput14 WD3[0] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput25 WD3[1] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
Xinput36 WD3[2] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
XFILLER_0_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput47 opcode[0] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_4
XFILLER_0_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold809 rf.registers\[20\]\[20\] VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7543__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5360__B1 _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5338__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5060_ rf.registers\[4\]\[18\] rf.registers\[5\]\[18\] rf.registers\[6\]\[18\] rf.registers\[7\]\[18\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__mux4_1
XANTENNA__6683__A _3230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8374__S _4132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8750_ clknet_leaf_29_clk _0934_ VGND VGND VPWR VPWR rf.registers\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_5962_ _2675_ _2703_ _2347_ VGND VGND VPWR VPWR _2704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7701_ _3025_ net779 _3808_ VGND VGND VPWR VPWR _3810_ sky130_fd_sc_hd__mux2_1
X_4913_ _1668_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__clkbuf_4
X_8681_ clknet_leaf_64_clk _0865_ VGND VGND VPWR VPWR rf.registers\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5893_ net114 _1542_ _1558_ VGND VGND VPWR VPWR _2638_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7632_ _3773_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_43_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6622__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4844_ _1205_ _1599_ _1057_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5274__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7563_ _3019_ net470 _3736_ VGND VGND VPWR VPWR _3737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4775_ rf.registers\[28\]\[9\] rf.registers\[29\]\[9\] rf.registers\[30\]\[9\] rf.registers\[31\]\[9\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__mux4_2
XFILLER_0_43_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9302_ clknet_leaf_24_clk _0462_ VGND VGND VPWR VPWR rf.registers\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6514_ net634 _3103_ _3157_ VGND VGND VPWR VPWR _3163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7494_ _3699_ VGND VGND VPWR VPWR _3700_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_151_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9233_ clknet_leaf_30_clk _0393_ VGND VGND VPWR VPWR rf.registers\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_151_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6445_ net152 _3118_ _3114_ VGND VGND VPWR VPWR _3119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9164_ clknet_leaf_45_clk _0324_ VGND VGND VPWR VPWR rf.registers\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6376_ net29 VGND VGND VPWR VPWR _3071_ sky130_fd_sc_hd__clkbuf_2
X_8115_ _4029_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5327_ _2064_ _2082_ VGND VGND VPWR VPWR _2083_ sky130_fd_sc_hd__and2_1
XANTENNA__5329__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9095_ clknet_leaf_66_clk _0255_ VGND VGND VPWR VPWR rf.registers\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_8046_ net432 _3462_ _3989_ VGND VGND VPWR VPWR _3993_ sky130_fd_sc_hd__mux2_1
X_5258_ _1766_ _2013_ _1672_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_71_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5189_ rf.registers\[24\]\[28\] rf.registers\[25\]\[28\] rf.registers\[26\]\[28\]
+ rf.registers\[27\]\[28\] _1882_ _1884_ VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_3_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6603__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8948_ clknet_leaf_30_clk _0108_ VGND VGND VPWR VPWR rf.registers\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5501__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5002__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire82 _1667_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
X_8879_ clknet_leaf_10_clk _0039_ VGND VGND VPWR VPWR rf.registers\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5265__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1_A _1181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4560__B _1315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5590__B1 _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4987__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7363__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4288__A _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8194__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5847__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6442__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5256__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5058__S _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _1299_ _1315_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4897__S net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4491_ rf.registers\[8\]\[20\] rf.registers\[9\]\[20\] rf.registers\[10\]\[20\] rf.registers\[11\]\[20\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__mux4_1
Xhold606 rf.registers\[17\]\[26\] VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5559__S1 _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold617 rf.registers\[27\]\[12\] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold628 rf.registers\[28\]\[8\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 rf.registers\[27\]\[25\] VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6230_ _2955_ _2503_ _2956_ VGND VGND VPWR VPWR _2957_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6161_ _2015_ _2889_ VGND VGND VPWR VPWR _2892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5112_ _1866_ _1867_ _1713_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__mux2_1
X_6092_ _2812_ _2817_ _2808_ VGND VGND VPWR VPWR _2827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5043_ _1167_ VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8802_ clknet_leaf_55_clk _0986_ VGND VGND VPWR VPWR rf.registers\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6994_ net263 _3103_ _3413_ VGND VGND VPWR VPWR _3419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4298__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8733_ clknet_leaf_14_clk _0917_ VGND VGND VPWR VPWR rf.registers\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5945_ _2684_ _2686_ _2160_ VGND VGND VPWR VPWR _2688_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7448__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5757__A _2305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6352__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8664_ clknet_leaf_11_clk _0848_ VGND VGND VPWR VPWR rf.registers\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5876_ _1839_ _2211_ _2248_ VGND VGND VPWR VPWR _2622_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5247__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7615_ _3075_ net1001 _3758_ VGND VGND VPWR VPWR _3764_ sky130_fd_sc_hd__mux2_1
X_4827_ rf.registers\[4\]\[16\] rf.registers\[5\]\[16\] rf.registers\[6\]\[16\] rf.registers\[7\]\[16\]
+ net1158 _1183_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__mux4_1
X_8595_ clknet_leaf_35_clk _0779_ VGND VGND VPWR VPWR rf.registers\[22\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xclone28 _1637_ VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7546_ _3727_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
X_4758_ rf.registers\[16\]\[8\] rf.registers\[17\]\[8\] rf.registers\[18\]\[8\] rf.registers\[19\]\[8\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__mux4_2
XFILLER_0_133_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4470__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8279__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7477_ _3073_ net1032 _3686_ VGND VGND VPWR VPWR _3691_ sky130_fd_sc_hd__mux2_1
XANTENNA__5492__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7183__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4689_ _1439_ _1441_ _1444_ _1254_ _1170_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9216_ clknet_leaf_69_clk _0376_ VGND VGND VPWR VPWR rf.registers\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6428_ net43 VGND VGND VPWR VPWR _3107_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5875__B2 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9147_ clknet_leaf_36_clk _0307_ VGND VGND VPWR VPWR rf.registers\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6359_ _3059_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7911__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9078_ clknet_leaf_33_clk _0238_ VGND VGND VPWR VPWR rf.registers\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6527__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8029_ _3011_ net679 _3974_ VGND VGND VPWR VPWR _3983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4289__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clone45_A _1219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5667__A _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4571__A _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_73_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7093__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4510__S _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5410__S0 _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5866__B2 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7821__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5577__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7268__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5730_ _2080_ _2448_ VGND VGND VPWR VPWR _2483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5229__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5661_ _2332_ _2415_ VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__xnor2_1
X_7400_ _3627_ VGND VGND VPWR VPWR _3650_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4612_ _1366_ _1367_ _1199_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__mux2_1
X_8380_ net429 _3454_ _4169_ VGND VGND VPWR VPWR _4170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5592_ _1146_ VGND VGND VPWR VPWR _2347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7331_ _3590_ VGND VGND VPWR VPWR _3613_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4543_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__inv_2
Xhold403 rf.registers\[8\]\[26\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold414 rf.registers\[13\]\[23\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold425 rf.registers\[7\]\[25\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold436 rf.registers\[30\]\[10\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
X_7262_ _3576_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4474_ _1189_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__and2_1
Xhold447 rf.registers\[12\]\[18\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5401__S0 _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9001_ clknet_leaf_50_clk _0161_ VGND VGND VPWR VPWR rf.registers\[31\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold458 rf.registers\[2\]\[17\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 rf.registers\[27\]\[0\] VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _2934_ _2940_ VGND VGND VPWR VPWR _2941_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7193_ _3516_ VGND VGND VPWR VPWR _3539_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _2033_ _2874_ VGND VGND VPWR VPWR _2876_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_5_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8128__A _4024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6075_ _1838_ _2783_ VGND VGND VPWR VPWR _2811_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _1733_ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__8562__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6034__A1 _1874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6034__B2 _1858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6977_ net413 _3015_ _3375_ VGND VGND VPWR VPWR _3409_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8716_ clknet_leaf_45_clk _0900_ VGND VGND VPWR VPWR rf.registers\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5928_ _2428_ _2288_ VGND VGND VPWR VPWR _2672_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_66_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8647_ clknet_leaf_5_clk _0831_ VGND VGND VPWR VPWR rf.registers\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5859_ _2404_ _2605_ _2591_ _2356_ VGND VGND VPWR VPWR _2606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6810__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8578_ clknet_leaf_58_clk _0762_ VGND VGND VPWR VPWR rf.registers\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7529_ _3718_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold970 rf.registers\[2\]\[24\] VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7641__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold981 rf.registers\[23\]\[29\] VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 rf.registers\[28\]\[24\] VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4520__A1 _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5459__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5397__A _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4587__A1 _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4682__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6720__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6956__A _3375_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7551__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5860__A _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7787__A _3843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6900_ _3368_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8382__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7880_ _3904_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_74_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6831_ net399 _3145_ _3326_ VGND VGND VPWR VPWR _3332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9550_ clknet_leaf_28_clk _0710_ VGND VGND VPWR VPWR rf.registers\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4578__A1 _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6762_ _3075_ net748 _3289_ VGND VGND VPWR VPWR _3295_ sky130_fd_sc_hd__mux2_1
X_8501_ _4233_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5713_ _2255_ _2463_ _2465_ _2373_ VGND VGND VPWR VPWR _2466_ sky130_fd_sc_hd__o211a_1
X_9481_ clknet_leaf_51_clk _0641_ VGND VGND VPWR VPWR rf.registers\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6693_ _3258_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7726__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6630__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8432_ net774 _3508_ _4191_ VGND VGND VPWR VPWR _4197_ sky130_fd_sc_hd__mux2_1
X_5644_ _1842_ _1838_ _1799_ VGND VGND VPWR VPWR _2399_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5754__B _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8363_ _4160_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__clkbuf_1
X_5575_ _1669_ _1660_ VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__or2_2
XANTENNA__5246__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold200 rf.registers\[7\]\[5\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold211 rf.registers\[3\]\[5\] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
X_7314_ _3604_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4526_ _1280_ _1281_ _1198_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__mux2_1
Xhold222 rf.registers\[7\]\[31\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
X_8294_ _3143_ net901 _4119_ VGND VGND VPWR VPWR _4124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold233 rf.registers\[0\]\[2\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold244 rf.registers\[24\]\[9\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 rf.registers\[5\]\[24\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
X_7245_ _3046_ net426 _3566_ VGND VGND VPWR VPWR _3568_ sky130_fd_sc_hd__mux2_1
X_4457_ _1038_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__clkbuf_8
Xhold266 rf.registers\[6\]\[15\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold277 rf.registers\[7\]\[28\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5770__A _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold288 rf.registers\[11\]\[16\] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 rf.registers\[1\]\[15\] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7176_ _3530_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
X_4388_ _1025_ _1135_ _1139_ _1143_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6127_ _2719_ _2731_ VGND VGND VPWR VPWR _2860_ sky130_fd_sc_hd__and2_1
X_6058_ _2373_ _2476_ _2789_ _2794_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_68_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8292__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5009_ _1761_ _1764_ _1697_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4361__S0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4325__S _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5010__A _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4664__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5156__S _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7371__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4296__A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7400__A _3627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5839__B _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4655__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4407__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5360_ _1685_ _2115_ _1696_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4311_ rf.registers\[28\]\[5\] rf.registers\[29\]\[5\] rf.registers\[30\]\[5\] rf.registers\[31\]\[5\]
+ net101 _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5291_ rf.registers\[24\]\[3\] rf.registers\[25\]\[3\] rf.registers\[26\]\[3\] rf.registers\[27\]\[3\]
+ _1674_ _1691_ VGND VGND VPWR VPWR _2047_ sky130_fd_sc_hd__mux4_1
XANTENNA__6485__A1 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7030_ net343 _3139_ _3435_ VGND VGND VPWR VPWR _3438_ sky130_fd_sc_hd__mux2_1
X_8981_ clknet_leaf_35_clk _0141_ VGND VGND VPWR VPWR rf.registers\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_143_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4343__S0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7932_ net482 _3485_ _3927_ VGND VGND VPWR VPWR _3932_ sky130_fd_sc_hd__mux2_1
XANTENNA__4934__A _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7310__A _3590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7863_ _3895_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6814_ net418 _3128_ _3315_ VGND VGND VPWR VPWR _3323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7794_ net156 _3483_ _3855_ VGND VGND VPWR VPWR _3859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9533_ clknet_leaf_15_clk _0693_ VGND VGND VPWR VPWR rf.registers\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6745_ _3058_ net1041 _3278_ VGND VGND VPWR VPWR _3286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7456__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5765__A _2323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9464_ clknet_leaf_21_clk _0624_ VGND VGND VPWR VPWR rf.registers\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6676_ _3249_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8415_ net520 _3491_ _4180_ VGND VGND VPWR VPWR _4188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5627_ _2378_ _2381_ _1877_ VGND VGND VPWR VPWR _2382_ sky130_fd_sc_hd__mux2_1
X_9395_ clknet_leaf_35_clk _0555_ VGND VGND VPWR VPWR rf.registers\[24\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5071__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4723__A1 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8346_ _4151_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5558_ _2310_ _2313_ net4 VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4509_ _1261_ _1264_ _1259_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__mux2_1
X_8277_ _3126_ net1068 _4108_ VGND VGND VPWR VPWR _4115_ sky130_fd_sc_hd__mux2_1
X_5489_ _1697_ _2240_ _2242_ _2244_ _1729_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__a221o_1
XANTENNA__7191__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7228_ _3029_ net271 _3555_ VGND VGND VPWR VPWR _3559_ sky130_fd_sc_hd__mux2_1
X_7159_ _3521_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4582__S0 _1267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6535__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4637__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5675__A _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8197__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6219__A1 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6445__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5978__A0 _2650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4860_ _1614_ _1615_ _1189_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__8392__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4791_ rf.registers\[24\]\[10\] rf.registers\[25\]\[10\] rf.registers\[26\]\[10\]
+ rf.registers\[27\]\[10\] _1041_ _1043_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_31_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5585__A _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7276__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6530_ _3171_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6180__S _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6461_ _3129_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8200_ _4074_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5053__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5412_ rf.registers\[12\]\[12\] rf.registers\[13\]\[12\] rf.registers\[14\]\[12\]
+ rf.registers\[15\]\[12\] _2117_ _2118_ VGND VGND VPWR VPWR _2168_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9180_ clknet_leaf_18_clk _0340_ VGND VGND VPWR VPWR rf.registers\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6392_ _3081_ net613 _3065_ VGND VGND VPWR VPWR _3082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8131_ net1143 _3479_ _4036_ VGND VGND VPWR VPWR _4038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5343_ _1167_ _2098_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__or2_1
XANTENNA__4929__A _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5524__S _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8062_ _4001_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__clkbuf_1
X_5274_ rf.registers\[0\]\[24\] rf.registers\[1\]\[24\] rf.registers\[2\]\[24\] rf.registers\[3\]\[24\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__mux4_1
X_7013_ net237 _3122_ _3424_ VGND VGND VPWR VPWR _3429_ sky130_fd_sc_hd__mux2_1
XANTENNA__4564__S0 _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6355__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8964_ clknet_leaf_47_clk _0124_ VGND VGND VPWR VPWR rf.registers\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7915_ net478 _3468_ _3916_ VGND VGND VPWR VPWR _3923_ sky130_fd_sc_hd__mux2_1
X_8895_ clknet_leaf_71_clk _0055_ VGND VGND VPWR VPWR rf.registers\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7846_ _3886_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4619__S1 _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5197__A1 _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7777_ net341 _3466_ _3844_ VGND VGND VPWR VPWR _3850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4989_ _1686_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4603__S _1214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6728_ _3041_ net772 _3267_ VGND VGND VPWR VPWR _3277_ sky130_fd_sc_hd__mux2_1
X_9516_ clknet_leaf_45_clk _0676_ VGND VGND VPWR VPWR rf.registers\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9447_ clknet_leaf_5_clk _0607_ VGND VGND VPWR VPWR rf.registers\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6659_ _3240_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9378_ clknet_leaf_59_clk _0538_ VGND VGND VPWR VPWR rf.registers\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5942__B _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8329_ _4142_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4555__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7949__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4307__S0 _1026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4858__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7096__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5609__S _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8126__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput15 WD3[10] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xinput26 WD3[20] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput37 WD3[30] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xinput48 opcode[1] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_4
XFILLER_0_109_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5360__A1 _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4794__S0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5344__S _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5961_ _2161_ _2142_ VGND VGND VPWR VPWR _2703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7700_ _3809_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8390__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4912_ net82 VGND VGND VPWR VPWR _1668_ sky130_fd_sc_hd__buf_2
XANTENNA__6903__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8680_ clknet_leaf_63_clk _0864_ VGND VGND VPWR VPWR rf.registers\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5892_ _2627_ _2629_ _2637_ _2621_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__o22a_1
XFILLER_0_75_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7631_ net924 _3454_ _3772_ VGND VGND VPWR VPWR _3773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4843_ _1597_ _1598_ _1036_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5274__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4423__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7562_ _3735_ VGND VGND VPWR VPWR _3736_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__6204__A _1958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4774_ rf.registers\[16\]\[9\] rf.registers\[17\]\[9\] rf.registers\[18\]\[9\] rf.registers\[19\]\[9\]
+ net106 _1073_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__mux4_2
XFILLER_0_28_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9301_ clknet_leaf_34_clk _0461_ VGND VGND VPWR VPWR rf.registers\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6513_ _3162_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7493_ _3193_ _3626_ VGND VGND VPWR VPWR _3699_ sky130_fd_sc_hd__nand2_4
XFILLER_0_71_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7734__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9232_ clknet_leaf_12_clk _0392_ VGND VGND VPWR VPWR rf.registers\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6444_ net17 VGND VGND VPWR VPWR _3118_ sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_9_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9163_ clknet_leaf_4_clk _0323_ VGND VGND VPWR VPWR rf.registers\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6375_ _3070_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8114_ net648 _3462_ _4025_ VGND VGND VPWR VPWR _4029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5326_ _1168_ _2081_ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__nand2_1
X_9094_ clknet_leaf_0_clk _0254_ VGND VGND VPWR VPWR rf.registers\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8045_ _3992_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__clkbuf_1
X_5257_ _2011_ _2012_ _1745_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5188_ _1800_ _1943_ VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8947_ clknet_leaf_33_clk _0107_ VGND VGND VPWR VPWR rf.registers\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7909__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8878_ clknet_leaf_41_clk _0038_ VGND VGND VPWR VPWR rf.registers\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8356__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7829_ net193 _3450_ _3843_ VGND VGND VPWR VPWR _3877_ sky130_fd_sc_hd__mux2_1
XANTENNA__5515__A1_N _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5265__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_rebuffer18_A _1464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4569__A _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4776__S0 _1290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8475__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4528__S0 net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4302__C1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5802__C1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7819__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4700__S0 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4724__A1_N _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5847__B _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5339__S net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5256__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6024__A _1858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7858__A0 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4490_ _1242_ _1245_ _1187_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__mux2_2
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold607 rf.registers\[23\]\[20\] VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold618 rf.registers\[14\]\[27\] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 rf.registers\[16\]\[30\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6160_ _2890_ VGND VGND VPWR VPWR _2891_ sky130_fd_sc_hd__inv_2
XANTENNA__4541__C1 _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7086__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5111_ rf.registers\[12\]\[16\] rf.registers\[13\]\[16\] rf.registers\[14\]\[16\]
+ rf.registers\[15\]\[16\] _1720_ _1723_ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__mux4_1
XANTENNA__8283__A0 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6091_ _2528_ _2823_ _2731_ _2824_ _2825_ VGND VGND VPWR VPWR _2826_ sky130_fd_sc_hd__a221o_1
X_5042_ _1729_ _1789_ _1797_ VGND VGND VPWR VPWR _1798_ sky130_fd_sc_hd__a21oi_2
XANTENNA__5192__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4844__B1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5103__A _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8801_ clknet_leaf_56_clk _0985_ VGND VGND VPWR VPWR rf.registers\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6597__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6993_ _3418_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5944_ _2686_ _2684_ _2160_ VGND VGND VPWR VPWR _2687_ sky130_fd_sc_hd__and3_1
X_8732_ clknet_leaf_17_clk _0916_ VGND VGND VPWR VPWR rf.registers\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6349__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8663_ clknet_leaf_24_clk _0847_ VGND VGND VPWR VPWR rf.registers\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5875_ _2607_ _2614_ _2620_ _2621_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__o22a_1
XANTENNA__5249__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5247__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7614_ _3763_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4826_ _1213_ _1581_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8594_ clknet_leaf_38_clk _0778_ VGND VGND VPWR VPWR rf.registers\[22\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xclone18 _1089_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone29 _1200_ VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7545_ _3073_ net781 _3722_ VGND VGND VPWR VPWR _3727_ sky130_fd_sc_hd__mux2_1
X_4757_ rf.registers\[20\]\[8\] rf.registers\[21\]\[8\] rf.registers\[22\]\[8\] rf.registers\[23\]\[8\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__mux4_2
XANTENNA__7464__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7849__A0 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7476_ _3690_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
X_4688_ _1442_ _1443_ _1211_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__mux2_1
XANTENNA__8510__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9215_ clknet_leaf_70_clk _0375_ VGND VGND VPWR VPWR rf.registers\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5324__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6427_ _3106_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4758__S0 _1026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4389__A _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9146_ clknet_leaf_37_clk _0306_ VGND VGND VPWR VPWR rf.registers\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6358_ _3058_ net322 _3044_ VGND VGND VPWR VPWR _3059_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7077__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5309_ rf.registers\[20\]\[2\] rf.registers\[21\]\[2\] rf.registers\[22\]\[2\] rf.registers\[23\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__mux4_1
XANTENNA__6808__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9077_ clknet_leaf_42_clk _0237_ VGND VGND VPWR VPWR rf.registers\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6289_ net34 VGND VGND VPWR VPWR _3011_ sky130_fd_sc_hd__clkbuf_4
X_8028_ _3982_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5183__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7639__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6543__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clone38_A _1065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5454__A1_N _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5159__S _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6760__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4771__C1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5410__S1 _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8265__A0 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6718__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5174__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7549__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5858__A _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5229__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5660_ _2413_ _2414_ VGND VGND VPWR VPWR _2415_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4611_ rf.registers\[0\]\[25\] rf.registers\[1\]\[25\] rf.registers\[2\]\[25\] rf.registers\[3\]\[25\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5591_ _2344_ _2345_ VGND VGND VPWR VPWR _2346_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7284__S _3554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7330_ _3612_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
X_4542_ _1286_ _1170_ _1297_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__a21o_4
XFILLER_0_52_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold404 rf.registers\[15\]\[20\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 rf.registers\[1\]\[24\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
X_7261_ _3062_ net625 _3566_ VGND VGND VPWR VPWR _3576_ sky130_fd_sc_hd__mux2_1
Xhold426 rf.registers\[18\]\[11\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ rf.registers\[4\]\[28\] rf.registers\[5\]\[28\] rf.registers\[6\]\[28\] rf.registers\[7\]\[28\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__mux4_1
Xhold437 rf.registers\[20\]\[12\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 rf.registers\[31\]\[4\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9000_ clknet_leaf_46_clk _0160_ VGND VGND VPWR VPWR rf.registers\[31\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold459 rf.registers\[18\]\[4\] VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _2885_ _2936_ _2939_ VGND VGND VPWR VPWR _2940_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5401__S1 _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7192_ _3538_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8256__A0 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6143_ _2033_ _2874_ VGND VGND VPWR VPWR _2875_ sky130_fd_sc_hd__nor2_1
XANTENNA__6628__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4937__A _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6806__A1 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _1838_ _2783_ _2768_ _1820_ VGND VGND VPWR VPWR _2810_ sky130_fd_sc_hd__a211o_1
X_5025_ _1168_ _1780_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_146_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6976_ _3408_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8715_ clknet_leaf_5_clk _0899_ VGND VGND VPWR VPWR rf.registers\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5927_ _2669_ _2670_ VGND VGND VPWR VPWR _2671_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8646_ clknet_leaf_1_clk _0830_ VGND VGND VPWR VPWR rf.registers\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_5858_ _1111_ _2102_ VGND VGND VPWR VPWR _2605_ sky130_fd_sc_hd__nor2_2
XFILLER_0_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4809_ rf.registers\[12\]\[11\] rf.registers\[13\]\[11\] rf.registers\[14\]\[11\]
+ rf.registers\[15\]\[11\] _1052_ _1053_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7194__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8577_ clknet_leaf_58_clk _0761_ VGND VGND VPWR VPWR rf.registers\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5789_ _2271_ _2538_ VGND VGND VPWR VPWR _2539_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5707__S _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7528_ _3056_ net975 _3711_ VGND VGND VPWR VPWR _3718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7459_ _3681_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold960 rf.registers\[25\]\[23\] VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 rf.registers\[22\]\[10\] VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 rf.registers\[22\]\[24\] VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 rf.registers\[22\]\[11\] VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__dlygate4sd3_1
X_9129_ clknet_leaf_50_clk _0289_ VGND VGND VPWR VPWR rf.registers\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_110_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7369__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5459__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6273__S _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6733__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output76_A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6448__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5472__B1 _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4492__A _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6830_ _3331_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6761_ _3294_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5712_ _1148_ _2368_ _2369_ _2464_ _2336_ VGND VGND VPWR VPWR _2465_ sky130_fd_sc_hd__a311o_1
X_8500_ net253 net31 _4227_ VGND VGND VPWR VPWR _4233_ sky130_fd_sc_hd__mux2_1
XANTENNA__6911__S _3339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9480_ clknet_leaf_52_clk _0640_ VGND VGND VPWR VPWR rf.registers\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6692_ net923 _3143_ _3253_ VGND VGND VPWR VPWR _3258_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_114_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5643_ _1842_ _1798_ net82 VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__o21a_1
X_8431_ _4196_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5754__C _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8362_ net749 _3506_ _4155_ VGND VGND VPWR VPWR _4160_ sky130_fd_sc_hd__mux2_1
X_5574_ _2041_ _1666_ _2103_ _2329_ VGND VGND VPWR VPWR _2330_ sky130_fd_sc_hd__o22a_1
X_7313_ _3046_ net966 _3602_ VGND VGND VPWR VPWR _3604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold201 rf.registers\[25\]\[3\] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4525_ rf.registers\[16\]\[26\] rf.registers\[17\]\[26\] rf.registers\[18\]\[26\]
+ rf.registers\[19\]\[26\] net1158 _1183_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__mux4_2
Xhold212 rf.registers\[20\]\[0\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
X_8293_ _4123_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold223 rf.registers\[1\]\[23\] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold234 rf.registers\[16\]\[22\] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold245 rf.registers\[16\]\[13\] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
X_7244_ _3567_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__9395__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold256 rf.registers\[13\]\[27\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _1209_ _1210_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__mux2_2
Xhold267 rf.registers\[10\]\[2\] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold278 rf.registers\[9\]\[19\] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold289 rf.registers\[24\]\[27\] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7175_ net140 _3479_ _3528_ VGND VGND VPWR VPWR _3530_ sky130_fd_sc_hd__mux2_1
XANTENNA__6358__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4387_ _1088_ _1142_ net8 VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_123_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6126_ _2791_ _2858_ _2501_ VGND VGND VPWR VPWR _2859_ sky130_fd_sc_hd__mux2_1
X_6057_ _2651_ _2731_ _2792_ _2496_ _2793_ VGND VGND VPWR VPWR _2794_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5008_ _1762_ _1763_ _1726_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4361__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5498__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7189__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7204__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5310__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6959_ net809 _3137_ _3398_ VGND VGND VPWR VPWR _3400_ sky130_fd_sc_hd__mux2_1
XANTENNA__7917__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6821__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8629_ clknet_leaf_35_clk _0813_ VGND VGND VPWR VPWR rf.registers\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4341__S _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6191__A1 _1996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7652__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_141_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7691__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold790 rf.registers\[8\]\[12\] VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5129__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8483__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7099__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7827__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6731__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6182__A1 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4310_ A2[1] VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5290_ rf.registers\[28\]\[3\] rf.registers\[29\]\[3\] rf.registers\[30\]\[3\] rf.registers\[31\]\[3\]
+ _1674_ _1691_ VGND VGND VPWR VPWR _2046_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5693__B1 _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8980_ clknet_leaf_42_clk _0140_ VGND VGND VPWR VPWR rf.registers\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_143_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7931_ _3931_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4343__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7862_ _3120_ net691 _3891_ VGND VGND VPWR VPWR _3895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6813_ _3322_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7793_ _3858_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4950__A _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9532_ clknet_leaf_16_clk _0692_ VGND VGND VPWR VPWR rf.registers\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6744_ _3285_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6675_ net735 _3126_ _3242_ VGND VGND VPWR VPWR _3249_ sky130_fd_sc_hd__mux2_1
X_9463_ clknet_leaf_23_clk _0623_ VGND VGND VPWR VPWR rf.registers\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5257__S _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7038__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8414_ _4187_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__clkbuf_1
X_5626_ _2379_ _2380_ VGND VGND VPWR VPWR _2381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9394_ clknet_leaf_39_clk _0554_ VGND VGND VPWR VPWR rf.registers\[24\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5557_ _2311_ _2312_ _1684_ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8345_ net412 _3489_ _4144_ VGND VGND VPWR VPWR _4151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4508_ rf.registers\[24\]\[21\] rf.registers\[25\]\[21\] rf.registers\[26\]\[21\]
+ rf.registers\[27\]\[21\] _1262_ _1263_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__mux4_2
XANTENNA__5359__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8276_ _4114_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5488_ _1712_ _2243_ _1716_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__o21a_1
XANTENNA__7673__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7227_ _3558_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4397__A _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4439_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7158_ net386 _3462_ _3517_ VGND VGND VPWR VPWR _3521_ sky130_fd_sc_hd__mux2_1
XANTENNA__4582__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6109_ _2806_ _2841_ _2842_ VGND VGND VPWR VPWR _2843_ sky130_fd_sc_hd__a21oi_1
XANTENNA__6816__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7089_ _3455_ VGND VGND VPWR VPWR _3477_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__5436__B1 _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5021__A _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7647__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8332__A _4132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clone20_A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_rebuffer48_A _1217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7382__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7664__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6726__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5522__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7557__S _3699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4790_ rf.registers\[28\]\[10\] rf.registers\[29\]\[10\] rf.registers\[30\]\[10\]
+ rf.registers\[31\]\[10\] net93 _1043_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__mux4_2
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_18 _3194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6460_ net158 _3128_ _3114_ VGND VGND VPWR VPWR _3129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6155__B2 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5411_ rf.registers\[8\]\[12\] rf.registers\[9\]\[12\] rf.registers\[10\]\[12\] rf.registers\[11\]\[12\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2167_ sky130_fd_sc_hd__mux4_1
XANTENNA__8388__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6391_ net34 VGND VGND VPWR VPWR _3081_ sky130_fd_sc_hd__buf_2
XANTENNA__7292__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8130_ _4037_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5342_ _1638_ _2097_ VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8061_ net581 _3476_ _4000_ VGND VGND VPWR VPWR _4001_ sky130_fd_sc_hd__mux2_1
X_5273_ rf.registers\[4\]\[24\] rf.registers\[5\]\[24\] rf.registers\[6\]\[24\] rf.registers\[7\]\[24\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__mux4_1
X_7012_ _3428_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6636__S _3194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4945__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5540__S _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5418__B1 _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8963_ clknet_leaf_66_clk _0123_ VGND VGND VPWR VPWR rf.registers\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7914_ _3922_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__clkbuf_1
X_8894_ clknet_leaf_0_clk _0054_ VGND VGND VPWR VPWR rf.registers\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7845_ _3103_ net859 _3880_ VGND VGND VPWR VPWR _3886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6371__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7776_ _3849_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__clkbuf_1
X_4988_ _1740_ _1743_ _1697_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9515_ clknet_leaf_6_clk _0675_ VGND VGND VPWR VPWR rf.registers\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6727_ _3276_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7991__A _3951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9446_ clknet_leaf_72_clk _0606_ VGND VGND VPWR VPWR rf.registers\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6658_ net435 _3109_ _3231_ VGND VGND VPWR VPWR _3240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8298__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5609_ _2359_ _2362_ _2363_ VGND VGND VPWR VPWR _2364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9377_ clknet_leaf_58_clk _0537_ VGND VGND VPWR VPWR rf.registers\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6589_ _3203_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8328_ net687 _3472_ _4133_ VGND VGND VPWR VPWR _4142_ sky130_fd_sc_hd__mux2_1
XANTENNA__6400__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8259_ _4105_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7930__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5016__A _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5657__B1 _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4555__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6546__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4855__A _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8800__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8071__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4307__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5504__S0 _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7377__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4491__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput16 WD3[11] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XANTENNA__6137__A1 _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput27 WD3[21] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 WD3[31] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4794__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4765__A _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5960_ _2421_ _2690_ _2691_ _2695_ _2702_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__o32a_1
X_4911_ _1171_ _1153_ _1157_ _1161_ _1165_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__a32oi_4
X_5891_ _2633_ _2636_ VGND VGND VPWR VPWR _2637_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7630_ _3771_ VGND VGND VPWR VPWR _3772_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4842_ rf.registers\[0\]\[17\] rf.registers\[1\]\[17\] rf.registers\[2\]\[17\] rf.registers\[3\]\[17\]
+ net1158 _1183_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4387__B1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4773_ rf.registers\[20\]\[9\] rf.registers\[21\]\[9\] rf.registers\[22\]\[9\] rf.registers\[23\]\[9\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__mux4_2
X_7561_ _3155_ _3553_ VGND VGND VPWR VPWR _3735_ sky130_fd_sc_hd__nand2b_4
XTAP_TAPCELL_ROW_138_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9300_ clknet_leaf_42_clk _0460_ VGND VGND VPWR VPWR rf.registers\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6512_ net362 _3101_ _3157_ VGND VGND VPWR VPWR _3162_ sky130_fd_sc_hd__mux2_1
XANTENNA__6128__A1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7492_ _3698_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9231_ clknet_leaf_27_clk _0391_ VGND VGND VPWR VPWR rf.registers\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6443_ _3117_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_151_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9162_ clknet_leaf_7_clk _0322_ VGND VGND VPWR VPWR rf.registers\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6374_ _3069_ net1120 _3065_ VGND VGND VPWR VPWR _3070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8113_ _4028_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__clkbuf_1
X_5325_ net1163 _2080_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__nor2_1
X_9093_ clknet_leaf_57_clk _0253_ VGND VGND VPWR VPWR rf.registers\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8044_ net1037 _3460_ _3989_ VGND VGND VPWR VPWR _3992_ sky130_fd_sc_hd__mux2_1
X_5256_ rf.registers\[0\]\[25\] rf.registers\[1\]\[25\] rf.registers\[2\]\[25\] rf.registers\[3\]\[25\]
+ _1767_ _1768_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5187_ net1163 _1942_ VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__and2b_1
XANTENNA__4862__A1 _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7800__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8946_ clknet_leaf_25_clk _0106_ VGND VGND VPWR VPWR rf.registers\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8877_ clknet_leaf_41_clk _0037_ VGND VGND VPWR VPWR rf.registers\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7828_ _3876_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7759_ _3083_ net1133 _3830_ VGND VGND VPWR VPWR _3840_ sky130_fd_sc_hd__mux2_1
XANTENNA__4473__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5590__A2 _2160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__9479__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9429_ clknet_leaf_32_clk _0589_ VGND VGND VPWR VPWR rf.registers\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5445__S _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4776__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7660__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4528__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4585__A _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4700__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6305__A _3022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7555__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7835__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold608 rf.registers\[28\]\[1\] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold619 rf.registers\[10\]\[6\] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5110_ rf.registers\[8\]\[16\] rf.registers\[9\]\[16\] rf.registers\[10\]\[16\] rf.registers\[11\]\[16\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__mux4_1
X_6090_ _2102_ _2523_ VGND VGND VPWR VPWR _2825_ sky130_fd_sc_hd__nor2_1
X_5041_ _1791_ _1793_ _1796_ _1697_ _1671_ VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_53_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4844__A1 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5192__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8800_ clknet_leaf_68_clk _0984_ VGND VGND VPWR VPWR rf.registers\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5103__B _1858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6992_ net638 _3101_ _3413_ VGND VGND VPWR VPWR _3418_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4831__A1_N _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8731_ clknet_leaf_22_clk _0915_ VGND VGND VPWR VPWR rf.registers\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_5943_ _2536_ _2657_ _2685_ _2683_ VGND VGND VPWR VPWR _2686_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8662_ clknet_leaf_33_clk _0846_ VGND VGND VPWR VPWR rf.registers\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_5874_ _2333_ VGND VGND VPWR VPWR _2621_ sky130_fd_sc_hd__buf_4
XFILLER_0_118_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7613_ _3073_ net1074 _3758_ VGND VGND VPWR VPWR _3763_ sky130_fd_sc_hd__mux2_1
X_4825_ _1579_ _1580_ _1287_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__mux2_1
X_8593_ clknet_leaf_41_clk _0777_ VGND VGND VPWR VPWR rf.registers\[22\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7745__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclone19 A2[0] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_16
X_7544_ _3726_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4756_ _1495_ _1511_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__and2_4
XFILLER_0_71_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4687_ rf.registers\[0\]\[22\] rf.registers\[1\]\[22\] rf.registers\[2\]\[22\] rf.registers\[3\]\[22\]
+ net132 _1175_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__mux4_1
X_7475_ _3071_ net1042 _3686_ VGND VGND VPWR VPWR _3690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9214_ clknet_leaf_71_clk _0374_ VGND VGND VPWR VPWR rf.registers\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6426_ net314 _3105_ _3093_ VGND VGND VPWR VPWR _3106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4758__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9145_ clknet_leaf_19_clk _0305_ VGND VGND VPWR VPWR rf.registers\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6357_ net22 VGND VGND VPWR VPWR _3058_ sky130_fd_sc_hd__clkbuf_2
X_5308_ _1167_ _2063_ VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__or2_1
X_9076_ clknet_leaf_42_clk _0236_ VGND VGND VPWR VPWR rf.registers\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6288_ _3010_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__clkbuf_1
X_8027_ _3009_ net1139 _3974_ VGND VGND VPWR VPWR _3982_ sky130_fd_sc_hd__mux2_1
X_5239_ _1773_ _1990_ _1992_ _1994_ _1672_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__o221a_1
XANTENNA__5183__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8929_ clknet_leaf_56_clk _0089_ VGND VGND VPWR VPWR rf.registers\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4694__S0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7537__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6512__A1 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7390__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4519__S _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5174__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5204__A _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload3_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5858__B _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7528__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7565__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5874__A _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4610_ rf.registers\[4\]\[25\] rf.registers\[5\]\[25\] rf.registers\[6\]\[25\] rf.registers\[7\]\[25\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__mux4_1
X_5590_ _2144_ _2160_ _1668_ VGND VGND VPWR VPWR _2345_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4541_ _1289_ _1293_ _1296_ _1205_ _1025_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold405 rf.registers\[0\]\[26\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
X_7260_ _3575_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
X_4472_ _1224_ _1227_ _1187_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__mux2_4
XFILLER_0_123_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold416 rf.registers\[19\]\[23\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold427 rf.registers\[17\]\[24\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_36_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold438 rf.registers\[12\]\[17\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 rf.registers\[17\]\[25\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9024__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6211_ _2891_ _2937_ _2935_ _2938_ _2916_ VGND VGND VPWR VPWR _2939_ sky130_fd_sc_hd__o311a_1
XANTENNA__8396__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7191_ net892 _3495_ _3528_ VGND VGND VPWR VPWR _3538_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6909__S _3339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6142_ _1384_ _2873_ VGND VGND VPWR VPWR _2874_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_5_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _2769_ _2784_ VGND VGND VPWR VPWR _2809_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5024_ _1758_ _1779_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_146_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5490__A1 _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6019__B1 _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6644__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6975_ net502 _3013_ _3398_ VGND VGND VPWR VPWR _3408_ sky130_fd_sc_hd__mux2_1
XANTENNA__4676__S0 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8714_ clknet_leaf_8_clk _0898_ VGND VGND VPWR VPWR rf.registers\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5926_ _2663_ _2668_ VGND VGND VPWR VPWR _2670_ sky130_fd_sc_hd__nand2_1
XANTENNA__6990__A1 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8645_ clknet_leaf_53_clk _0829_ VGND VGND VPWR VPWR rf.registers\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5857_ _2390_ _2590_ VGND VGND VPWR VPWR _2604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7475__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4808_ rf.registers\[8\]\[11\] rf.registers\[9\]\[11\] rf.registers\[10\]\[11\] rf.registers\[11\]\[11\]
+ net117 _1053_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__mux4_1
X_8576_ clknet_leaf_69_clk _0760_ VGND VGND VPWR VPWR rf.registers\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5788_ net119 _2537_ VGND VGND VPWR VPWR _2538_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7527_ _3717_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
X_4739_ _1464_ _1480_ _1494_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7458_ _3054_ net670 _3675_ VGND VGND VPWR VPWR _3681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6409_ _3094_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__clkbuf_1
Xhold950 rf.registers\[25\]\[24\] VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 rf.registers\[30\]\[3\] VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__dlygate4sd3_1
X_7389_ _3644_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4600__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5723__S _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold972 rf.registers\[17\]\[23\] VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__dlygate4sd3_1
X_9128_ clknet_leaf_46_clk _0288_ VGND VGND VPWR VPWR rf.registers\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold983 rf.registers\[15\]\[19\] VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 rf.registers\[31\]\[16\] VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__dlygate4sd3_1
X_9059_ clknet_leaf_68_clk _0219_ VGND VGND VPWR VPWR rf.registers\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_110_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6554__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clone50_A _1172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4667__S0 net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5633__S _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output69_A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5472__A1 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7749__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6760_ _3073_ net653 _3289_ VGND VGND VPWR VPWR _3294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5711_ _2178_ _2362_ VGND VGND VPWR VPWR _2464_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6691_ _3257_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__clkbuf_1
X_8430_ net675 _3506_ _4191_ VGND VGND VPWR VPWR _4196_ sky130_fd_sc_hd__mux2_1
X_5642_ _2393_ _2396_ _1146_ VGND VGND VPWR VPWR _2397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8361_ _4159_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5754__D _1166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5573_ _2105_ _2253_ _2255_ _2328_ VGND VGND VPWR VPWR _2329_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_103_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7312_ _3603_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8477__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4524_ rf.registers\[20\]\[26\] rf.registers\[21\]\[26\] rf.registers\[22\]\[26\]
+ rf.registers\[23\]\[26\] net1156 _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__mux4_2
Xhold202 rf.registers\[5\]\[28\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
X_8292_ _3141_ net496 _4119_ VGND VGND VPWR VPWR _4123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold213 rf.registers\[7\]\[16\] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 rf.registers\[7\]\[29\] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 rf.registers\[20\]\[27\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 rf.registers\[21\]\[7\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
X_7243_ _3043_ net949 _3566_ VGND VGND VPWR VPWR _3567_ sky130_fd_sc_hd__mux2_1
XANTENNA__4948__A _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4455_ _1198_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5543__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold257 rf.registers\[2\]\[18\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4499__C1 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold268 rf.registers\[24\]\[8\] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 rf.registers\[2\]\[10\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4386_ _1140_ _1141_ _1107_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7174_ _3529_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6125_ _2820_ _2857_ _1147_ VGND VGND VPWR VPWR _2858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6056_ _2458_ _2738_ VGND VGND VPWR VPWR _2793_ sky130_fd_sc_hd__nor2_1
XANTENNA__5779__A _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6374__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5007_ rf.registers\[24\]\[21\] rf.registers\[25\]\[21\] rf.registers\[26\]\[21\]
+ rf.registers\[27\]\[21\] _1676_ _1681_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__mux4_1
XANTENNA__4683__A _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8401__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5498__B _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6958_ _3399_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5310__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5909_ _2468_ _2530_ _2475_ _2503_ VGND VGND VPWR VPWR _2654_ sky130_fd_sc_hd__a31o_1
XANTENNA__4974__B1 _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6889_ net617 _3134_ _3362_ VGND VGND VPWR VPWR _3363_ sky130_fd_sc_hd__mux2_1
XANTENNA__5718__S _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4622__S _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8628_ clknet_leaf_38_clk _0812_ VGND VGND VPWR VPWR rf.registers\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6403__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5074__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8559_ _4263_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4821__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5377__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold780 rf.registers\[4\]\[11\] VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 rf.registers\[21\]\[18\] VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7979__A0 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5129__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4888__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6284__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4593__A _1334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6954__A1 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8004__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6167__C1 _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7843__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4812__S0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5693__A1 _1145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6983__A _3412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_143_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7930_ net164 _3483_ _3927_ VGND VGND VPWR VPWR _3931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7861_ _3894_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7198__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6812_ net794 _3126_ _3315_ VGND VGND VPWR VPWR _3322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7792_ net147 _3481_ _3855_ VGND VGND VPWR VPWR _3858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9531_ clknet_leaf_21_clk _0691_ VGND VGND VPWR VPWR rf.registers\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6743_ _3056_ net1151 _3278_ VGND VGND VPWR VPWR _3285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9462_ clknet_leaf_24_clk _0622_ VGND VGND VPWR VPWR rf.registers\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6674_ _3248_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5056__S0 _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8413_ net895 _3489_ _4180_ VGND VGND VPWR VPWR _4187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5625_ _1167_ _1943_ VGND VGND VPWR VPWR _2380_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9393_ clknet_leaf_40_clk _0553_ VGND VGND VPWR VPWR rf.registers\[24\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4803__S0 _1072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7753__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8344_ _4150_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__clkbuf_1
X_5556_ rf.registers\[24\]\[5\] rf.registers\[25\]\[5\] rf.registers\[26\]\[5\] rf.registers\[27\]\[5\]
+ _1702_ _1678_ VGND VGND VPWR VPWR _2312_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4507_ _1221_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8275_ _3124_ net1109 _4108_ VGND VGND VPWR VPWR _4114_ sky130_fd_sc_hd__mux2_1
X_5487_ rf.registers\[0\]\[9\] rf.registers\[1\]\[9\] rf.registers\[2\]\[9\] rf.registers\[3\]\[9\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__mux4_1
XANTENNA__5359__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7226_ _3027_ net988 _3555_ VGND VGND VPWR VPWR _3558_ sky130_fd_sc_hd__mux2_1
X_4438_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7157_ _3520_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4369_ _1024_ _1116_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__o21ai_4
X_6108_ _1779_ _2829_ VGND VGND VPWR VPWR _2842_ sky130_fd_sc_hd__and2b_1
X_7088_ net15 VGND VGND VPWR VPWR _3476_ sky130_fd_sc_hd__buf_2
XANTENNA__5436__A1 _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6039_ _1669_ _1821_ _1860_ VGND VGND VPWR VPWR _2777_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer50 net1169 VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__7189__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7928__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6936__A1 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5448__S _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4352__S _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6133__A _2038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clone13_A _1181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8494__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6624__A0 _3073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6308__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5522__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6927__A1 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5286__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 _3375_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5038__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7573__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5410_ _2162_ _2163_ _2164_ _2165_ _1711_ _1716_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6390_ _3080_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ _1640_ _2088_ _2096_ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__o21ai_4
XANTENNA_clkbuf_leaf_71_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4498__A _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5093__S _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8060_ _3988_ VGND VGND VPWR VPWR _4000_ sky130_fd_sc_hd__clkbuf_8
X_5272_ _1901_ _2027_ _1717_ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__a21o_1
XANTENNA__5210__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5666__A1 _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7011_ net364 _3120_ _3424_ VGND VGND VPWR VPWR _3428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6917__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5418__A1 _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8962_ clknet_leaf_59_clk _0122_ VGND VGND VPWR VPWR rf.registers\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8602__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7913_ net456 _3466_ _3916_ VGND VGND VPWR VPWR _3922_ sky130_fd_sc_hd__mux2_1
X_8893_ clknet_leaf_14_clk _0053_ VGND VGND VPWR VPWR rf.registers\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6652__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7844_ _3885_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4961__A _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7775_ net180 _3464_ _3844_ VGND VGND VPWR VPWR _3849_ sky130_fd_sc_hd__mux2_1
XANTENNA__5268__S _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4987_ _1741_ _1742_ _1739_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9514_ clknet_leaf_8_clk _0674_ VGND VGND VPWR VPWR rf.registers\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6726_ _3039_ net684 _3267_ VGND VGND VPWR VPWR _3276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9445_ clknet_leaf_61_clk _0605_ VGND VGND VPWR VPWR rf.registers\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6657_ _3239_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6888__A _3339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7483__S _3686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5608_ _1877_ VGND VGND VPWR VPWR _2363_ sky130_fd_sc_hd__buf_4
X_9376_ clknet_leaf_60_clk _0536_ VGND VGND VPWR VPWR rf.registers\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6588_ _3037_ net987 _3195_ VGND VGND VPWR VPWR _3203_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_39_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8327_ _4141_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__clkbuf_1
X_5539_ _2293_ _2294_ _2044_ VGND VGND VPWR VPWR _2295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8258_ _3107_ net782 _4097_ VGND VGND VPWR VPWR _4105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7209_ _3547_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6827__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8189_ _4068_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5504__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7658__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6562__S _3179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4491__S1 _1203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput17 WD3[12] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5906__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput28 WD3[22] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
Xinput39 WD3[3] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XANTENNA__4810__S _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5440__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5896__A1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5222__A1_N _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6737__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output51_A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6038__A _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4910_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__buf_2
X_5890_ _2598_ _2618_ _2617_ _2635_ VGND VGND VPWR VPWR _2636_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4841_ rf.registers\[4\]\[17\] rf.registers\[5\]\[17\] rf.registers\[6\]\[17\] rf.registers\[7\]\[17\]
+ net1158 _1183_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4387__A1 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7560_ _3734_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4772_ _1519_ _1025_ _1527_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__o21a_4
XFILLER_0_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6511_ _3161_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7491_ _3087_ net459 _3663_ VGND VGND VPWR VPWR _3698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9230_ clknet_leaf_29_clk _0390_ VGND VGND VPWR VPWR rf.registers\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5336__B1 _1655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6442_ net685 _3116_ _3114_ VGND VGND VPWR VPWR _3117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9161_ clknet_leaf_47_clk _0321_ VGND VGND VPWR VPWR rf.registers\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6373_ net28 VGND VGND VPWR VPWR _3069_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8112_ net825 _3460_ _4025_ VGND VGND VPWR VPWR _4028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5324_ net5 _2071_ _2079_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__a21oi_4
X_9092_ clknet_leaf_62_clk _0252_ VGND VGND VPWR VPWR rf.registers\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8043_ _3991_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4956__A _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5255_ rf.registers\[4\]\[25\] rf.registers\[5\]\[25\] rf.registers\[6\]\[25\] rf.registers\[7\]\[25\]
+ _1895_ _1897_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5186_ _1777_ _1933_ _1941_ VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7261__A0 _3062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8945_ clknet_leaf_44_clk _0105_ VGND VGND VPWR VPWR rf.registers\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4691__A _1430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8876_ clknet_leaf_49_clk _0036_ VGND VGND VPWR VPWR rf.registers\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7827_ net198 _3448_ _3866_ VGND VGND VPWR VPWR _3876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7758_ _3839_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4473__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6709_ _3266_ VGND VGND VPWR VPWR _3267_ sky130_fd_sc_hd__buf_4
X_7689_ net618 _3446_ _3794_ VGND VGND VPWR VPWR _3803_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9428_ clknet_leaf_29_clk _0588_ VGND VGND VPWR VPWR rf.registers\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8102__S _3988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9359_ clknet_leaf_10_clk _0519_ VGND VGND VPWR VPWR rf.registers\[20\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7242__A _3554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4302__B2 _1038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7388__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5802__A1 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5566__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4540__S _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold609 rf.registers\[23\]\[13\] VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7851__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4541__B2 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5371__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5040_ _1794_ _1795_ _1739_ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7243__A0 _3043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6991_ _3417_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7298__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8730_ clknet_leaf_17_clk _0914_ VGND VGND VPWR VPWR rf.registers\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4715__S _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5942_ _1464_ _2411_ VGND VGND VPWR VPWR _2685_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8661_ clknet_leaf_32_clk _0845_ VGND VGND VPWR VPWR rf.registers\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5873_ _2617_ _2619_ VGND VGND VPWR VPWR _2620_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7612_ _3762_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4824_ rf.registers\[12\]\[16\] rf.registers\[13\]\[16\] rf.registers\[14\]\[16\]
+ rf.registers\[15\]\[16\] _1191_ _1174_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8592_ clknet_leaf_14_clk _0776_ VGND VGND VPWR VPWR rf.registers\[22\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7543_ _3071_ net979 _3722_ VGND VGND VPWR VPWR _3726_ sky130_fd_sc_hd__mux2_1
X_4755_ _1239_ _1502_ _1506_ _1510_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_145_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7474_ _3689_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
X_4686_ rf.registers\[4\]\[22\] rf.registers\[5\]\[22\] rf.registers\[6\]\[22\] rf.registers\[7\]\[22\]
+ net132 _1175_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9213_ clknet_leaf_3_clk _0373_ VGND VGND VPWR VPWR rf.registers\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6425_ net42 VGND VGND VPWR VPWR _3105_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7761__S _3807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9144_ clknet_leaf_11_clk _0304_ VGND VGND VPWR VPWR rf.registers\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6356_ _3057_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__clkbuf_1
X_5307_ _1638_ _2062_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__or2_1
XANTENNA__6377__S _3065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9075_ clknet_leaf_35_clk _0235_ VGND VGND VPWR VPWR rf.registers\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6287_ net186 _3009_ _3007_ VGND VGND VPWR VPWR _3010_ sky130_fd_sc_hd__mux2_1
X_8026_ _3981_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__clkbuf_1
X_5238_ _1901_ _1993_ _1766_ VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__a21o_1
X_5169_ _1169_ _1924_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7785__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8928_ clknet_leaf_69_clk _0088_ VGND VGND VPWR VPWR rf.registers\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4694__S1 _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8859_ clknet_leaf_22_clk _0019_ VGND VGND VPWR VPWR rf.registers\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7936__S _3927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5548__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6141__A _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4771__B2 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6287__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4596__A _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6276__B2 _2472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6028__B2 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5787__B1 _2536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6200__A1 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4540_ _1294_ _1295_ _1287_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold406 rf.registers\[1\]\[16\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
X_4471_ _1225_ _1226_ _1178_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__mux2_1
Xhold417 rf.registers\[11\]\[2\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7581__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold428 rf.registers\[22\]\[4\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold439 rf.registers\[11\]\[9\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6210_ _1996_ _2903_ _2917_ VGND VGND VPWR VPWR _2938_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7190_ _3537_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6141_ _2595_ _2872_ VGND VGND VPWR VPWR _2873_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_5_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7464__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6072_ _2806_ _2807_ VGND VGND VPWR VPWR _2808_ sky130_fd_sc_hd__or2_1
X_5023_ _1672_ _1765_ _1772_ _1778_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__6925__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4373__S0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6019__A1 _1127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6974_ _3407_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4676__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8713_ clknet_leaf_65_clk _0897_ VGND VGND VPWR VPWR rf.registers\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_5925_ _2663_ _2668_ VGND VGND VPWR VPWR _2669_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4450__B1 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6660__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8644_ clknet_leaf_51_clk _0828_ VGND VGND VPWR VPWR rf.registers\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5856_ _2587_ _2589_ _2592_ _2603_ _2408_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__o32a_1
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4807_ _1559_ _1560_ _1561_ _1562_ _1048_ _1050_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__mux4_2
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8575_ clknet_leaf_73_clk _0759_ VGND VGND VPWR VPWR rf.registers\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5787_ net95 net131 _2536_ VGND VGND VPWR VPWR _2537_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7526_ _3054_ net727 _3711_ VGND VGND VPWR VPWR _3717_ sky130_fd_sc_hd__mux2_1
X_4738_ _1215_ _1485_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7457_ _3680_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__clkbuf_1
X_4669_ _1214_ _1424_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7491__S _3663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6408_ net681 _3089_ _3093_ VGND VGND VPWR VPWR _3094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold940 rf.registers\[21\]\[25\] VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__dlygate4sd3_1
X_7388_ _3052_ net503 _3639_ VGND VGND VPWR VPWR _3644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold951 rf.registers\[20\]\[9\] VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 rf.registers\[24\]\[19\] VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4600__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9127_ clknet_leaf_66_clk _0287_ VGND VGND VPWR VPWR rf.registers\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold973 rf.registers\[22\]\[25\] VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ net16 VGND VGND VPWR VPWR _3046_ sky130_fd_sc_hd__buf_2
Xhold984 rf.registers\[14\]\[15\] VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 rf.registers\[30\]\[27\] VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__dlygate4sd3_1
X_9058_ clknet_leaf_59_clk _0218_ VGND VGND VPWR VPWR rf.registers\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_110_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5024__B _1779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8009_ _3972_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6835__S _3326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4667__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7666__S _3783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5941__B1 _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4845__A1_N _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6745__S _3278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_128_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5710_ _2354_ _2359_ _2178_ VGND VGND VPWR VPWR _2463_ sky130_fd_sc_hd__mux2_1
X_6690_ net450 _3141_ _3253_ VGND VGND VPWR VPWR _3257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5641_ _2394_ _2395_ VGND VGND VPWR VPWR _2396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7921__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5096__S _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8360_ net712 _3504_ _4155_ VGND VGND VPWR VPWR _4159_ sky130_fd_sc_hd__mux2_1
X_5572_ _2289_ _2326_ _2327_ VGND VGND VPWR VPWR _2328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7311_ _3043_ net818 _3602_ VGND VGND VPWR VPWR _3603_ sky130_fd_sc_hd__mux2_1
X_4523_ _1073_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8291_ _4122_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold203 rf.registers\[19\]\[24\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 rf.registers\[2\]\[5\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold225 rf.registers\[5\]\[27\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
X_7242_ _3554_ VGND VGND VPWR VPWR _3566_ sky130_fd_sc_hd__buf_4
Xhold236 rf.registers\[8\]\[30\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ rf.registers\[0\]\[29\] rf.registers\[1\]\[29\] rf.registers\[2\]\[29\] rf.registers\[3\]\[29\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold247 rf.registers\[3\]\[23\] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 rf.registers\[15\]\[17\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 rf.registers\[6\]\[27\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7173_ net298 _3476_ _3528_ VGND VGND VPWR VPWR _3529_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4385_ rf.registers\[0\]\[1\] rf.registers\[1\]\[1\] rf.registers\[2\]\[1\] rf.registers\[3\]\[1\]
+ net102 _1090_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5125__A _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6124_ _2394_ _2392_ VGND VGND VPWR VPWR _2857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6055_ _2718_ _2791_ _2501_ VGND VGND VPWR VPWR _2792_ sky130_fd_sc_hd__mux2_1
XANTENNA__4964__A _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5999__B1 _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6660__A1 _3111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5006_ rf.registers\[28\]\[21\] rf.registers\[29\]\[21\] rf.registers\[30\]\[21\]
+ rf.registers\[31\]\[21\] _1676_ _1681_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_68_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6957_ net702 _3134_ _3398_ VGND VGND VPWR VPWR _3399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5908_ _1087_ _2652_ VGND VGND VPWR VPWR _2653_ sky130_fd_sc_hd__and2_1
XANTENNA__4974__A1 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6888_ _3339_ VGND VGND VPWR VPWR _3362_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5839_ _2335_ _2586_ VGND VGND VPWR VPWR _2587_ sky130_fd_sc_hd__nor2_1
X_8627_ clknet_leaf_36_clk _0811_ VGND VGND VPWR VPWR rf.registers\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5074__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7218__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8558_ net755 net27 _4255_ VGND VGND VPWR VPWR _4263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4821__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7509_ _3037_ net505 _3700_ VGND VGND VPWR VPWR _3708_ sky130_fd_sc_hd__mux2_1
X_8489_ _4204_ VGND VGND VPWR VPWR _4227_ sky130_fd_sc_hd__buf_4
XANTENNA__5734__S _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7515__A _3699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8110__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold770 rf.registers\[12\]\[22\] VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 rf.registers\[20\]\[19\] VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 rf.registers\[28\]\[2\] VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5035__A _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4888__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7600__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7396__S _3639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8081__A _3988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8156__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4812__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7419__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7860_ _3118_ net1050 _3891_ VGND VGND VPWR VPWR _3894_ sky130_fd_sc_hd__mux2_1
X_6811_ _3321_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__clkbuf_1
X_7791_ _3857_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5819__S _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6742_ _3284_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__clkbuf_1
X_9530_ clknet_leaf_18_clk _0690_ VGND VGND VPWR VPWR rf.registers\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8147__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9461_ clknet_leaf_31_clk _0621_ VGND VGND VPWR VPWR rf.registers\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6673_ net997 _3124_ _3242_ VGND VGND VPWR VPWR _3248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5056__S1 _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8412_ _4186_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__clkbuf_1
X_5624_ _1799_ _1924_ VGND VGND VPWR VPWR _2379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9392_ clknet_leaf_4_clk _0552_ VGND VGND VPWR VPWR rf.registers\[24\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4803__S1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8343_ net816 _3487_ _4144_ VGND VGND VPWR VPWR _4150_ sky130_fd_sc_hd__mux2_1
X_5555_ rf.registers\[28\]\[5\] rf.registers\[29\]\[5\] rf.registers\[30\]\[5\] rf.registers\[31\]\[5\]
+ _2050_ _1678_ VGND VGND VPWR VPWR _2311_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4959__A _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5554__S _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4506_ _1219_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__buf_12
X_8274_ _4113_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5486_ _1739_ _2241_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__or2_1
X_7225_ _3557_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_4437_ _1066_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7156_ net400 _3460_ _3517_ VGND VGND VPWR VPWR _3520_ sky130_fd_sc_hd__mux2_1
X_4368_ _1118_ _1120_ _1123_ _1037_ net8 VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a221o_1
X_6107_ _2829_ _1779_ VGND VGND VPWR VPWR _2841_ sky130_fd_sc_hd__or2b_1
XANTENNA__4319__S0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7087_ _3475_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
X_4299_ rf.registers\[12\]\[4\] rf.registers\[13\]\[4\] rf.registers\[14\]\[4\] rf.registers\[15\]\[4\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__mux4_1
XANTENNA__7070__A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6038_ _2102_ _2445_ VGND VGND VPWR VPWR _2776_ sky130_fd_sc_hd__nor2_1
Xrebuffer40 net121 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer51 _1277_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7989_ _3111_ net927 _3952_ VGND VGND VPWR VPWR _3962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5464__S _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4730__S0 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5286__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8015__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8129__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5038__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4779__A _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5374__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5340_ _2090_ _2092_ _2095_ net4 net5 VGND VGND VPWR VPWR _2096_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5271_ rf.registers\[8\]\[24\] rf.registers\[9\]\[24\] rf.registers\[10\]\[24\] rf.registers\[11\]\[24\]
+ _1881_ _1883_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__mux4_1
X_7010_ _3427_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5210__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4718__S _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8961_ clknet_leaf_57_clk _0121_ VGND VGND VPWR VPWR rf.registers\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7912_ _3921_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6933__S _3376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4721__S0 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8892_ clknet_leaf_16_clk _0052_ VGND VGND VPWR VPWR rf.registers\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_90_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7843_ _3101_ net243 _3880_ VGND VGND VPWR VPWR _3885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7774_ _3848_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4986_ rf.registers\[24\]\[22\] rf.registers\[25\]\[22\] rf.registers\[26\]\[22\]
+ rf.registers\[27\]\[22\] _1734_ _1735_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9513_ clknet_leaf_63_clk _0673_ VGND VGND VPWR VPWR rf.registers\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6725_ _3275_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7879__A0 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6656_ net356 _3107_ _3231_ VGND VGND VPWR VPWR _3239_ sky130_fd_sc_hd__mux2_1
X_9444_ clknet_leaf_62_clk _0604_ VGND VGND VPWR VPWR rf.registers\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5607_ _2360_ _2361_ VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__and2_1
X_9375_ clknet_leaf_73_clk _0535_ VGND VGND VPWR VPWR rf.registers\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6587_ _3202_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4788__S0 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8326_ net763 _3470_ _4133_ VGND VGND VPWR VPWR _4141_ sky130_fd_sc_hd__mux2_1
X_5538_ rf.registers\[24\]\[4\] rf.registers\[25\]\[4\] rf.registers\[26\]\[4\] rf.registers\[27\]\[4\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2294_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_76_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8257_ _4104_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5469_ rf.registers\[4\]\[8\] rf.registers\[5\]\[8\] rf.registers\[6\]\[8\] rf.registers\[7\]\[8\]
+ _1734_ _1735_ VGND VGND VPWR VPWR _2225_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5657__A2 _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7208_ net275 _3444_ _3539_ VGND VGND VPWR VPWR _3547_ sky130_fd_sc_hd__mux2_1
X_8188_ net179 _3468_ _4061_ VGND VGND VPWR VPWR _4068_ sky130_fd_sc_hd__mux2_1
X_7139_ _3510_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4614__A1_N _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6843__S _3303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4712__S0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6144__A _2033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8531__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 WD3[13] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_138_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput29 WD3[23] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5440__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5223__A _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7849__S _3880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4840_ _1213_ _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4771_ _1521_ _1523_ _1526_ _1050_ net8 VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__a221o_1
XANTENNA__5584__A1 _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7584__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6510_ net1010 _3099_ _3157_ VGND VGND VPWR VPWR _3161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5837__C_N _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7490_ _3697_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5336__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6441_ net16 VGND VGND VPWR VPWR _3116_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9160_ clknet_leaf_63_clk _0320_ VGND VGND VPWR VPWR rf.registers\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6372_ _3068_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8111_ _4027_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8286__A0 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5323_ _2073_ _2075_ _2078_ net4 _1640_ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9091_ clknet_leaf_67_clk _0251_ VGND VGND VPWR VPWR rf.registers\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8042_ net313 _3458_ _3989_ VGND VGND VPWR VPWR _3991_ sky130_fd_sc_hd__mux2_1
X_5254_ _1773_ _2009_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5185_ _1935_ _1937_ _1940_ _1773_ _1671_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_71_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5133__A _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7759__S _3830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6663__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4972__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8944_ clknet_leaf_12_clk _0104_ VGND VGND VPWR VPWR rf.registers\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5272__B1 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8875_ clknet_leaf_2_clk _0035_ VGND VGND VPWR VPWR rf.registers\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7013__A1 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7826_ _3875_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4969_ rf.registers\[0\]\[23\] rf.registers\[1\]\[23\] rf.registers\[2\]\[23\] rf.registers\[3\]\[23\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__mux4_1
X_7757_ _3081_ net945 _3830_ VGND VGND VPWR VPWR _3839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6708_ _3020_ _3192_ VGND VGND VPWR VPWR _3266_ sky130_fd_sc_hd__nand2_4
XFILLER_0_117_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7688_ _3802_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_22_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5912__A1_N _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9427_ clknet_leaf_32_clk _0587_ VGND VGND VPWR VPWR rf.registers\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6639_ _3229_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5308__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9358_ clknet_leaf_42_clk _0518_ VGND VGND VPWR VPWR rf.registers\[20\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8277__A0 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8309_ _4131_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__clkbuf_1
X_9289_ clknet_leaf_52_clk _0449_ VGND VGND VPWR VPWR rf.registers\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8029__A0 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5043__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_70_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5566__A1 _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5110__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_146_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6818__A1 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6049__A _1820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7579__S _3736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8264__A _4096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6990_ net194 _3099_ _3413_ VGND VGND VPWR VPWR _3417_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5941_ net1159 net90 _2411_ _2683_ VGND VGND VPWR VPWR _2684_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5872_ _2229_ _2597_ _2598_ _2618_ VGND VGND VPWR VPWR _2619_ sky130_fd_sc_hd__a2bb2o_1
X_8660_ clknet_leaf_30_clk _0844_ VGND VGND VPWR VPWR rf.registers\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4823_ rf.registers\[8\]\[16\] rf.registers\[9\]\[16\] rf.registers\[10\]\[16\] rf.registers\[11\]\[16\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__mux4_1
X_7611_ _3071_ net1029 _3758_ VGND VGND VPWR VPWR _3762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8591_ clknet_leaf_10_clk _0775_ VGND VGND VPWR VPWR rf.registers\[22\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8203__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4754_ _1254_ _1509_ _1170_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__a21oi_1
X_7542_ _3725_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7473_ _3069_ net1106 _3686_ VGND VGND VPWR VPWR _3689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4685_ _1199_ _1440_ _1213_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5128__A _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9212_ clknet_leaf_16_clk _0372_ VGND VGND VPWR VPWR rf.registers\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6424_ _3104_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6658__S _3231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6355_ _3056_ net1094 _3044_ VGND VGND VPWR VPWR _3057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9143_ clknet_leaf_34_clk _0303_ VGND VGND VPWR VPWR rf.registers\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4967__A _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5306_ _1729_ _2049_ _2057_ _2061_ VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__o2bb2a_1
X_9074_ clknet_leaf_39_clk _0234_ VGND VGND VPWR VPWR rf.registers\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6286_ net33 VGND VGND VPWR VPWR _3009_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5237_ rf.registers\[0\]\[26\] rf.registers\[1\]\[26\] rf.registers\[2\]\[26\] rf.registers\[3\]\[26\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__mux4_1
X_8025_ _3002_ net977 _3974_ VGND VGND VPWR VPWR _3981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5168_ _1639_ _1923_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__or2_1
XANTENNA__7489__S _3663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5099_ rf.registers\[0\]\[17\] rf.registers\[1\]\[17\] rf.registers\[2\]\[17\] rf.registers\[3\]\[17\]
+ _1822_ _1823_ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_104_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8927_ clknet_leaf_71_clk _0087_ VGND VGND VPWR VPWR rf.registers\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5796__A1 _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8858_ clknet_leaf_20_clk _0018_ VGND VGND VPWR VPWR rf.registers\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5548__A1 _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7809_ net354 _3497_ _3866_ VGND VGND VPWR VPWR _3867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8789_ clknet_leaf_32_clk _0973_ VGND VGND VPWR VPWR rf.registers\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4641__S _1040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6422__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6568__S _3156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6276__A2 _2737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5331__S0 _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8023__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6332__A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7862__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4470_ rf.registers\[24\]\[28\] rf.registers\[25\]\[28\] rf.registers\[26\]\[28\]
+ rf.registers\[27\]\[28\] _1220_ _1222_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__mux4_1
XANTENNA__5398__S0 _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold407 rf.registers\[5\]\[18\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 rf.registers\[24\]\[10\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 rf.registers\[7\]\[26\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5382__S _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6140_ _1447_ _2871_ VGND VGND VPWR VPWR _2872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6071_ _1798_ _2805_ VGND VGND VPWR VPWR _2807_ sky130_fd_sc_hd__and2_1
X_5022_ _1773_ _1776_ _1777_ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4373__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7102__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6973_ net830 _3011_ _3398_ VGND VGND VPWR VPWR _3407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8712_ clknet_leaf_63_clk _0896_ VGND VGND VPWR VPWR rf.registers\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5924_ _2602_ _2665_ _2667_ VGND VGND VPWR VPWR _2668_ sky130_fd_sc_hd__o21a_1
XANTENNA__4450__A1 _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8643_ clknet_leaf_54_clk _0827_ VGND VGND VPWR VPWR rf.registers\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_66_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5855_ _2598_ _2602_ VGND VGND VPWR VPWR _2603_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5557__S _1684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4806_ rf.registers\[20\]\[11\] rf.registers\[21\]\[11\] rf.registers\[22\]\[11\]
+ rf.registers\[23\]\[11\] _1072_ _1073_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__mux4_2
X_8574_ clknet_leaf_0_clk _0758_ VGND VGND VPWR VPWR rf.registers\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5786_ _2411_ VGND VGND VPWR VPWR _2536_ sky130_fd_sc_hd__buf_2
XFILLER_0_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7525_ _3716_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
X_4737_ _1487_ _1489_ _1492_ _1213_ _1057_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5389__S0 _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7456_ _3052_ net367 _3675_ VGND VGND VPWR VPWR _3680_ sky130_fd_sc_hd__mux2_1
X_4668_ _1422_ _1423_ _1190_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6407_ _3092_ VGND VGND VPWR VPWR _3093_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold930 rf.registers\[22\]\[23\] VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5292__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7387_ _3643_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
Xhold941 rf.registers\[4\]\[31\] VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _1353_ _1354_ _1199_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7073__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold952 rf.registers\[11\]\[31\] VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 rf.registers\[4\]\[27\] VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9126_ clknet_leaf_0_clk _0286_ VGND VGND VPWR VPWR rf.registers\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6338_ _3045_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__clkbuf_1
Xhold974 rf.registers\[14\]\[29\] VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold985 rf.registers\[30\]\[21\] VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold996 rf.registers\[22\]\[30\] VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__dlygate4sd3_1
X_9057_ clknet_leaf_58_clk _0217_ VGND VGND VPWR VPWR rf.registers\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6269_ _2992_ _2993_ VGND VGND VPWR VPWR _2994_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_110_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8008_ _3130_ net873 _3963_ VGND VGND VPWR VPWR _3972_ sky130_fd_sc_hd__mux2_1
XANTENNA__8108__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5313__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7947__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6851__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5975__B _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5467__S _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5991__A _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5552__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4546__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7382__A0 _3046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5640_ _1668_ _1780_ VGND VGND VPWR VPWR _2395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5571_ _1803_ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7592__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7310_ _3590_ VGND VGND VPWR VPWR _3602_ sky130_fd_sc_hd__buf_4
X_4522_ _1256_ _1277_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__nand2_1
X_8290_ _3139_ net909 _4119_ VGND VGND VPWR VPWR _4122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold204 rf.registers\[12\]\[10\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold215 rf.registers\[0\]\[8\] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
X_7241_ _3565_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
Xhold226 rf.registers\[10\]\[14\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ rf.registers\[4\]\[29\] rf.registers\[5\]\[29\] rf.registers\[6\]\[29\] rf.registers\[7\]\[29\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__mux4_1
Xhold237 rf.registers\[1\]\[4\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold248 rf.registers\[0\]\[1\] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4499__B2 _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold259 rf.registers\[9\]\[5\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7172_ _3516_ VGND VGND VPWR VPWR _3528_ sky130_fd_sc_hd__clkbuf_8
X_4384_ rf.registers\[4\]\[1\] rf.registers\[5\]\[1\] rf.registers\[6\]\[1\] rf.registers\[7\]\[1\]
+ net102 _1090_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_148_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6123_ _2854_ _2855_ VGND VGND VPWR VPWR _2856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6936__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6054_ _2752_ _2790_ _1147_ VGND VGND VPWR VPWR _2791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5005_ _1759_ _1760_ _1726_ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__mux2_1
XANTENNA__4456__S _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5141__A _1693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7767__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6671__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6956_ _3375_ VGND VGND VPWR VPWR _3398_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_81_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5907_ _2458_ _2487_ _2651_ _2530_ VGND VGND VPWR VPWR _2652_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_81_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6887_ _3361_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8626_ clknet_leaf_39_clk _0810_ VGND VGND VPWR VPWR rf.registers\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5838_ _2105_ _2584_ _2487_ _2585_ VGND VGND VPWR VPWR _2586_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_91_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8557_ _4262_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5769_ _2518_ _2519_ VGND VGND VPWR VPWR _2520_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_101_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7508_ _3707_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8488_ _4226_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7439_ _3035_ net1026 _3664_ VGND VGND VPWR VPWR _3671_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7007__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold760 rf.registers\[4\]\[4\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 rf.registers\[0\]\[15\] VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold782 rf.registers\[20\]\[24\] VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 rf.registers\[22\]\[12\] VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd3_1
X_9109_ clknet_leaf_30_clk _0269_ VGND VGND VPWR VPWR rf.registers\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5750__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5534__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7677__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6167__A1 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output74_A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6756__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8092__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6810_ net348 _3124_ _3315_ VGND VGND VPWR VPWR _3321_ sky130_fd_sc_hd__mux2_1
XANTENNA__6491__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7790_ net138 _3479_ _3855_ VGND VGND VPWR VPWR _3857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6741_ _3054_ net1066 _3278_ VGND VGND VPWR VPWR _3284_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9460_ clknet_leaf_30_clk _0620_ VGND VGND VPWR VPWR rf.registers\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6672_ _3247_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__clkbuf_1
X_8411_ net946 _3487_ _4180_ VGND VGND VPWR VPWR _4186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4708__A2 _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5366__C1 _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5623_ _2377_ VGND VGND VPWR VPWR _2378_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9391_ clknet_leaf_8_clk _0551_ VGND VGND VPWR VPWR rf.registers\[24\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5835__S _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8342_ _4149_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8211__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5554_ _2308_ _2309_ _1684_ VGND VGND VPWR VPWR _2310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4505_ rf.registers\[28\]\[21\] rf.registers\[29\]\[21\] rf.registers\[30\]\[21\]
+ rf.registers\[31\]\[21\] _1220_ _1222_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5485_ rf.registers\[4\]\[9\] rf.registers\[5\]\[9\] rf.registers\[6\]\[9\] rf.registers\[7\]\[9\]
+ _1734_ _1735_ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__mux4_1
X_8273_ _3122_ net1014 _4108_ VGND VGND VPWR VPWR _4113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7224_ _3025_ net632 _3555_ VGND VGND VPWR VPWR _3557_ sky130_fd_sc_hd__mux2_1
X_4436_ _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__buf_12
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7155_ _3519_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
X_4367_ _1121_ _1122_ _1047_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__mux2_1
XANTENNA__8447__A _4204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6106_ _2838_ _2839_ VGND VGND VPWR VPWR _2840_ sky130_fd_sc_hd__nand2_1
X_7086_ net717 _3474_ _3456_ VGND VGND VPWR VPWR _3475_ sky130_fd_sc_hd__mux2_1
XANTENNA__4319__S1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4298_ rf.registers\[8\]\[4\] rf.registers\[9\]\[4\] rf.registers\[10\]\[4\] rf.registers\[11\]\[4\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__mux4_1
X_6037_ _2769_ _2774_ VGND VGND VPWR VPWR _2775_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5841__B1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer30 _2633_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer41 _2725_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__7497__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer52 net133 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7594__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7988_ _3961_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__clkbuf_1
X_6939_ _3389_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8609_ clknet_leaf_56_clk _0793_ VGND VGND VPWR VPWR rf.registers\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9589_ clknet_leaf_32_clk _0749_ VGND VGND VPWR VPWR rf.registers\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7649__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold590 rf.registers\[23\]\[2\] VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4885__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6576__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5480__S _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5507__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4730__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7200__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8031__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7870__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5270_ _1889_ _2025_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__and2_1
X_8960_ clknet_leaf_59_clk _0120_ VGND VGND VPWR VPWR rf.registers\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_7911_ net541 _3464_ _3916_ VGND VGND VPWR VPWR _3921_ sky130_fd_sc_hd__mux2_1
XANTENNA__4721__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8891_ clknet_leaf_34_clk _0051_ VGND VGND VPWR VPWR rf.registers\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7842_ _3884_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7773_ net373 _3462_ _3844_ VGND VGND VPWR VPWR _3848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4985_ rf.registers\[28\]\[22\] rf.registers\[29\]\[22\] rf.registers\[30\]\[22\]
+ rf.registers\[31\]\[22\] _1734_ _1735_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4485__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9512_ clknet_leaf_63_clk _0672_ VGND VGND VPWR VPWR rf.registers\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6724_ _3037_ net661 _3267_ VGND VGND VPWR VPWR _3275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9443_ clknet_leaf_61_clk _0603_ VGND VGND VPWR VPWR rf.registers\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6655_ _3238_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5565__S _2044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5606_ net82 _2272_ VGND VGND VPWR VPWR _2361_ sky130_fd_sc_hd__nand2_1
X_9374_ clknet_leaf_0_clk _0534_ VGND VGND VPWR VPWR rf.registers\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4788__S1 _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6586_ _3035_ net829 _3195_ VGND VGND VPWR VPWR _3202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8325_ _4140_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__clkbuf_1
X_5537_ rf.registers\[28\]\[4\] rf.registers\[29\]\[4\] rf.registers\[30\]\[4\] rf.registers\[31\]\[4\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2293_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8256_ _3105_ net883 _4097_ VGND VGND VPWR VPWR _4104_ sky130_fd_sc_hd__mux2_1
X_5468_ _1697_ _2223_ VGND VGND VPWR VPWR _2224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7207_ _3546_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_4419_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__buf_4
X_8187_ _4067_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5399_ _1711_ _2154_ _1655_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7138_ net270 _3442_ _3498_ VGND VGND VPWR VPWR _3510_ sky130_fd_sc_hd__mux2_1
X_7069_ _3463_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4712__S1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8116__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6425__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5042__A1 _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7955__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7319__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_rebuffer46_A _1166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 WD3[14] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_150_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5223__B _1978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6335__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4467__S0 _1220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6781__A1 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4770_ _1524_ _1525_ _1035_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5893__B _1542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6440_ _3115_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6070__A _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6533__A1 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7730__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5741__C1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6371_ _3067_ net793 _3065_ VGND VGND VPWR VPWR _3068_ sky130_fd_sc_hd__mux2_1
X_8110_ net1017 _3458_ _4025_ VGND VGND VPWR VPWR _4027_ sky130_fd_sc_hd__mux2_1
X_5322_ _2076_ _2077_ _1684_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__mux2_1
X_9090_ clknet_leaf_59_clk _0250_ VGND VGND VPWR VPWR rf.registers\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8041_ _3990_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__clkbuf_1
X_5253_ _2007_ _2008_ _1713_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__mux2_1
XANTENNA__7105__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5414__A _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5184_ _1938_ _1939_ _1713_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6944__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8943_ clknet_leaf_28_clk _0103_ VGND VGND VPWR VPWR rf.registers\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5272__A1 _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8874_ clknet_leaf_64_clk _0034_ VGND VGND VPWR VPWR rf.registers\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4480__C1 _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7825_ net469 _3446_ _3866_ VGND VGND VPWR VPWR _3875_ sky130_fd_sc_hd__mux2_1
XANTENNA__7775__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7756_ _3838_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4968_ rf.registers\[4\]\[23\] rf.registers\[5\]\[23\] rf.registers\[6\]\[23\] rf.registers\[7\]\[23\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6707_ _3265_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7687_ net584 _3444_ _3794_ VGND VGND VPWR VPWR _3802_ sky130_fd_sc_hd__mux2_1
X_4899_ net4 VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7076__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9426_ clknet_leaf_27_clk _0586_ VGND VGND VPWR VPWR rf.registers\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_2__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6638_ _3087_ net1112 _3194_ VGND VGND VPWR VPWR _3229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9357_ clknet_leaf_40_clk _0517_ VGND VGND VPWR VPWR rf.registers\[20\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6569_ _3191_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4630__S0 _1219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8308_ _3017_ net302 _4096_ VGND VGND VPWR VPWR _4131_ sky130_fd_sc_hd__mux2_1
X_9288_ clknet_leaf_47_clk _0448_ VGND VGND VPWR VPWR rf.registers\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8239_ _4094_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7015__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4697__S0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7685__S _3794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5110__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5933__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4549__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5419__A1_N _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6764__S _3289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8440__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5940_ _1480_ VGND VGND VPWR VPWR _2683_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5871_ _2600_ _2601_ VGND VGND VPWR VPWR _2618_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7610_ _3761_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4822_ _1574_ _1575_ _1576_ _1577_ _1287_ _1078_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__mux4_1
X_8590_ clknet_leaf_42_clk _0774_ VGND VGND VPWR VPWR rf.registers\[22\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7541_ _3069_ net1091 _3722_ VGND VGND VPWR VPWR _3725_ sky130_fd_sc_hd__mux2_1
X_4753_ _1507_ _1508_ _1211_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6506__A1 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7472_ _3688_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
X_4684_ rf.registers\[12\]\[22\] rf.registers\[13\]\[22\] rf.registers\[14\]\[22\]
+ rf.registers\[15\]\[22\] _1192_ _1195_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__mux4_1
X_9211_ clknet_leaf_34_clk _0371_ VGND VGND VPWR VPWR rf.registers\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6423_ net473 _3103_ _3093_ VGND VGND VPWR VPWR _3104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9142_ clknet_leaf_33_clk _0302_ VGND VGND VPWR VPWR rf.registers\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6354_ net21 VGND VGND VPWR VPWR _3056_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_73_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4628__A1_N _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5305_ _1699_ _2060_ _1670_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__o21ai_1
X_9073_ clknet_leaf_40_clk _0233_ VGND VGND VPWR VPWR rf.registers\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6285_ _3008_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8024_ _3980_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__clkbuf_1
X_5236_ _1889_ _1991_ VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__and2_1
XANTENNA__5493__A1 _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4983__A _1738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5167_ _1777_ _1912_ _1916_ _1922_ VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__o2bb2a_2
X_5098_ rf.registers\[4\]\[17\] rf.registers\[5\]\[17\] rf.registers\[6\]\[17\] rf.registers\[7\]\[17\]
+ _1822_ _1823_ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_104_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4679__S0 _1182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8926_ clknet_leaf_0_clk _0086_ VGND VGND VPWR VPWR rf.registers\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8857_ clknet_leaf_23_clk _0017_ VGND VGND VPWR VPWR rf.registers\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7808_ _3843_ VGND VGND VPWR VPWR _3866_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8788_ clknet_leaf_30_clk _0972_ VGND VGND VPWR VPWR rf.registers\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7739_ _3829_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4851__S0 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8498__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9409_ clknet_leaf_56_clk _0569_ VGND VGND VPWR VPWR rf.registers\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6849__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7170__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5181__B1 _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6584__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8422__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5331__S1 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8304__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5095__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4842__S0 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5398__S1 _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold408 rf.registers\[19\]\[29\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold419 rf.registers\[6\]\[11\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6070_ _1798_ _2805_ VGND VGND VPWR VPWR _2806_ sky130_fd_sc_hd__nor2_1
X_5021_ _1729_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__6019__A3 _2737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8413__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6972_ _3406_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6975__A1 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8711_ clknet_leaf_66_clk _0895_ VGND VGND VPWR VPWR rf.registers\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5923_ _2645_ _2642_ net129 _2635_ _2666_ VGND VGND VPWR VPWR _2667_ sky130_fd_sc_hd__a221oi_2
XTAP_TAPCELL_ROW_24_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8642_ clknet_leaf_55_clk _0826_ VGND VGND VPWR VPWR rf.registers\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4742__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5854_ _2600_ _2601_ VGND VGND VPWR VPWR _2602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9365__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4805_ rf.registers\[16\]\[11\] rf.registers\[17\]\[11\] rf.registers\[18\]\[11\]
+ rf.registers\[19\]\[11\] _1072_ _1073_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__mux4_2
X_8573_ clknet_leaf_14_clk _0757_ VGND VGND VPWR VPWR rf.registers\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5785_ _1059_ _1083_ VGND VGND VPWR VPWR _2535_ sky130_fd_sc_hd__and2_4
XFILLER_0_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4833__S0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5139__A _1689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7524_ _3052_ net998 _3711_ VGND VGND VPWR VPWR _3716_ sky130_fd_sc_hd__mux2_1
X_4736_ _1490_ _1491_ _1287_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6669__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7455_ _3679_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4978__A _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4667_ rf.registers\[12\]\[23\] rf.registers\[13\]\[23\] rf.registers\[14\]\[23\]
+ rf.registers\[15\]\[23\] net1164 _1268_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__mux4_1
XANTENNA__5389__S1 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6406_ _3090_ _3091_ VGND VGND VPWR VPWR _3092_ sky130_fd_sc_hd__nor2_4
Xhold920 rf.registers\[19\]\[1\] VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7386_ _3050_ net474 _3639_ VGND VGND VPWR VPWR _3643_ sky130_fd_sc_hd__mux2_1
Xhold931 rf.registers\[28\]\[12\] VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4598_ rf.registers\[16\]\[25\] rf.registers\[17\]\[25\] rf.registers\[18\]\[25\]
+ rf.registers\[19\]\[25\] _1351_ _1352_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__mux4_1
Xhold942 rf.registers\[29\]\[16\] VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 rf.registers\[30\]\[4\] VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9125_ clknet_leaf_62_clk _0285_ VGND VGND VPWR VPWR rf.registers\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6337_ _3043_ net1053 _3044_ VGND VGND VPWR VPWR _3045_ sky130_fd_sc_hd__mux2_1
Xhold964 rf.registers\[30\]\[20\] VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold975 rf.registers\[0\]\[16\] VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 rf.registers\[13\]\[16\] VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 rf.registers\[31\]\[20\] VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__dlygate4sd3_1
X_9056_ clknet_leaf_60_clk _0216_ VGND VGND VPWR VPWR rf.registers\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6268_ _1334_ _1904_ VGND VGND VPWR VPWR _2993_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8007_ _3971_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5219_ rf.registers\[0\]\[27\] rf.registers\[1\]\[27\] rf.registers\[2\]\[27\] rf.registers\[3\]\[27\]
+ _1895_ _1897_ VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__mux4_1
X_6199_ _2475_ _2591_ _2652_ _2737_ _2927_ VGND VGND VPWR VPWR _2928_ sky130_fd_sc_hd__a221o_1
XANTENNA__5602__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5313__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8909_ clknet_leaf_44_clk _0069_ VGND VGND VPWR VPWR rf.registers\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8124__S _4025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clone29_A _1200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7963__S _3938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4824__S0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_37_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5457__A1 _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5552__S1 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6957__A1 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5068__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5570_ _2307_ _2325_ VGND VGND VPWR VPWR _2326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4521_ _1239_ _1266_ _1272_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__6489__S _3135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold205 rf.registers\[7\]\[30\] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7240_ _3041_ net1051 _3555_ VGND VGND VPWR VPWR _3565_ sky130_fd_sc_hd__mux2_1
Xhold216 rf.registers\[7\]\[10\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ _1174_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold227 rf.registers\[3\]\[30\] VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 rf.registers\[17\]\[8\] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold249 rf.registers\[17\]\[28\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7171_ _3527_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4383_ _1038_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7902__A _3915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6122_ _2840_ _2844_ _2838_ VGND VGND VPWR VPWR _2855_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6053_ _1800_ _1821_ _2399_ VGND VGND VPWR VPWR _2790_ sky130_fd_sc_hd__o21a_1
XANTENNA__8209__S _4072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5004_ rf.registers\[16\]\[21\] rf.registers\[17\]\[21\] rf.registers\[18\]\[21\]
+ rf.registers\[19\]\[21\] _1676_ _1681_ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_68_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6952__S _3387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6948__A1 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6955_ _3397_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5620__A1 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5906_ _2648_ _2650_ _2501_ VGND VGND VPWR VPWR _2651_ sky130_fd_sc_hd__mux2_1
XANTENNA__4472__S _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6886_ net379 _3132_ _3351_ VGND VGND VPWR VPWR _3361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8625_ clknet_leaf_39_clk _0809_ VGND VGND VPWR VPWR rf.registers\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5837_ _1758_ _2331_ _1148_ VGND VGND VPWR VPWR _2585_ sky130_fd_sc_hd__or3b_1
XANTENNA__7783__S _3844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4806__S0 _1072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8556_ net917 net26 _4255_ VGND VGND VPWR VPWR _4262_ sky130_fd_sc_hd__mux2_1
X_5768_ _2511_ _2512_ _2509_ VGND VGND VPWR VPWR _2519_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7507_ _3035_ net861 _3700_ VGND VGND VPWR VPWR _3707_ sky130_fd_sc_hd__mux2_1
X_4719_ _1213_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8487_ net822 net24 _4216_ VGND VGND VPWR VPWR _4226_ sky130_fd_sc_hd__mux2_1
X_5699_ _2449_ _2451_ VGND VGND VPWR VPWR _2453_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7438_ _3670_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold750 rf.registers\[26\]\[29\] VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd3_1
X_7369_ _3033_ net1020 _3628_ VGND VGND VPWR VPWR _3634_ sky130_fd_sc_hd__mux2_1
Xhold761 rf.registers\[22\]\[9\] VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 rf.registers\[9\]\[27\] VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold783 rf.registers\[25\]\[20\] VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd3_1
X_9108_ clknet_leaf_30_clk _0268_ VGND VGND VPWR VPWR rf.registers\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold794 rf.registers\[26\]\[24\] VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9039_ clknet_leaf_9_clk _0199_ VGND VGND VPWR VPWR rf.registers\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6428__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5534__S1 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7023__S _3424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5298__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4382__S _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7693__S _3771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5470__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output67_A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4557__S _1199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8029__S _3974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5242__A _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7868__S _3891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6772__S _3266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6740_ _3283_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6671_ net570 _3122_ _3242_ VGND VGND VPWR VPWR _3247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8410_ _4185_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5622_ _1168_ _1905_ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9390_ clknet_leaf_41_clk _0550_ VGND VGND VPWR VPWR rf.registers\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5461__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8341_ net704 _3485_ _4144_ VGND VGND VPWR VPWR _4149_ sky130_fd_sc_hd__mux2_1
XANTENNA__8304__A0 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5553_ rf.registers\[16\]\[5\] rf.registers\[17\]\[5\] rf.registers\[18\]\[5\] rf.registers\[19\]\[5\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2309_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7108__S _3477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6012__S _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4504_ _1257_ _1258_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__mux2_1
XANTENNA__4321__A _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8272_ _4112_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5484_ _2238_ _2239_ _1685_ VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__mux2_1
X_7223_ _3556_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4435_ _1072_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__buf_12
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7154_ net454 _3458_ _3517_ VGND VGND VPWR VPWR _3519_ sky130_fd_sc_hd__mux2_1
X_4366_ rf.registers\[12\]\[2\] rf.registers\[13\]\[2\] rf.registers\[14\]\[2\] rf.registers\[15\]\[2\]
+ net101 _1066_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6105_ _1754_ _2837_ VGND VGND VPWR VPWR _2839_ sky130_fd_sc_hd__or2_1
X_7085_ net45 VGND VGND VPWR VPWR _3474_ sky130_fd_sc_hd__buf_2
X_4297_ _1043_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__buf_4
X_6036_ _2749_ _2771_ _2773_ VGND VGND VPWR VPWR _2774_ sky130_fd_sc_hd__a21bo_1
Xrebuffer31 _2724_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer42 _2745_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlymetal6s2s_1
X_7987_ _3109_ net791 _3952_ VGND VGND VPWR VPWR _3961_ sky130_fd_sc_hd__mux2_1
XANTENNA__7079__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6938_ net862 _3116_ _3387_ VGND VGND VPWR VPWR _3389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6869_ _3352_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8608_ clknet_leaf_68_clk _0792_ VGND VGND VPWR VPWR rf.registers\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9588_ clknet_leaf_30_clk _0748_ VGND VGND VPWR VPWR rf.registers\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8539_ net585 net17 _4244_ VGND VGND VPWR VPWR _4253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6857__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold580 rf.registers\[18\]\[0\] VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold591 rf.registers\[23\]\[30\] VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6158__A _1370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5507__S1 _2114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7282__A0 _3083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5997__A _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__S _3195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8312__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5443__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5671__S _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5823__A1 _2472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7598__S _3747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5823__B2 _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7910_ _3920_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__clkbuf_1
X_8890_ clknet_leaf_37_clk _0050_ VGND VGND VPWR VPWR rf.registers\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4904__A1_N _1640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7841_ _3099_ net455 _3880_ VGND VGND VPWR VPWR _3884_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7772_ _3847_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4316__A _1041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4984_ _1736_ _1737_ _1739_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9511_ clknet_leaf_66_clk _0671_ VGND VGND VPWR VPWR rf.registers\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6723_ _3274_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4485__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9442_ clknet_leaf_60_clk _0602_ VGND VGND VPWR VPWR rf.registers\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6654_ net410 _3105_ _3231_ VGND VGND VPWR VPWR _3238_ sky130_fd_sc_hd__mux2_1
XANTENNA__8222__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5434__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5605_ _1668_ _2324_ VGND VGND VPWR VPWR _2360_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9373_ clknet_leaf_15_clk _0533_ VGND VGND VPWR VPWR rf.registers\[20\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6585_ _3201_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8324_ net953 _3468_ _4133_ VGND VGND VPWR VPWR _4140_ sky130_fd_sc_hd__mux2_1
X_5536_ _2290_ _2291_ _2044_ VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8255_ _4103_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6677__S _3242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5467_ _2221_ _2222_ _1712_ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7206_ net511 _3442_ _3539_ VGND VGND VPWR VPWR _3546_ sky130_fd_sc_hd__mux2_1
X_4418_ _1073_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__buf_4
X_8186_ net277 _3466_ _4061_ VGND VGND VPWR VPWR _4067_ sky130_fd_sc_hd__mux2_1
X_5398_ rf.registers\[0\]\[13\] rf.registers\[1\]\[13\] rf.registers\[2\]\[13\] rf.registers\[3\]\[13\]
+ _1702_ _1678_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__mux4_1
X_7137_ _3509_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
X_4349_ _1043_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7264__A0 _3064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7068_ net303 _3462_ _3456_ VGND VGND VPWR VPWR _3463_ sky130_fd_sc_hd__mux2_1
X_6019_ _1127_ _2524_ _2737_ _2503_ VGND VGND VPWR VPWR _2758_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_107_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5578__B1 _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6441__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5425__S0 _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7971__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6058__A1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7255__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4467__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7447__A _3663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8042__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6351__A net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_40_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__5416__S0 _1718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7881__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6370_ net27 VGND VGND VPWR VPWR _3067_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5321_ rf.registers\[0\]\[2\] rf.registers\[1\]\[2\] rf.registers\[2\]\[2\] rf.registers\[3\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6497__S _3092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8040_ net294 _3454_ _3989_ VGND VGND VPWR VPWR _3990_ sky130_fd_sc_hd__mux2_1
X_5252_ rf.registers\[12\]\[25\] rf.registers\[13\]\[25\] rf.registers\[14\]\[25\]
+ rf.registers\[15\]\[25\] _1895_ _1897_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__mux4_1
X_5183_ rf.registers\[12\]\[29\] rf.registers\[13\]\[29\] rf.registers\[14\]\[29\]
+ rf.registers\[15\]\[29\] _1767_ _1768_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4745__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8942_ clknet_leaf_29_clk _0102_ VGND VGND VPWR VPWR rf.registers\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7121__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8873_ clknet_leaf_52_clk _0033_ VGND VGND VPWR VPWR rf.registers\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4480__B1 _1205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7824_ _3874_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6221__A1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4967_ _1722_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__buf_4
X_7755_ _3079_ net1077 _3830_ VGND VGND VPWR VPWR _3838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6706_ net563 _3017_ _3230_ VGND VGND VPWR VPWR _3265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5980__B1 _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7686_ _3801_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
X_4898_ net4 _1653_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5407__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9425_ clknet_leaf_42_clk _0585_ VGND VGND VPWR VPWR rf.registers\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6637_ _3228_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9356_ clknet_leaf_50_clk _0516_ VGND VGND VPWR VPWR rf.registers\[20\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6568_ net803 _3017_ _3156_ VGND VGND VPWR VPWR _3191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4630__S1 _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5519_ rf.registers\[16\]\[7\] rf.registers\[17\]\[7\] rf.registers\[18\]\[7\] rf.registers\[19\]\[7\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__mux4_1
X_8307_ _4130_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__clkbuf_1
X_9287_ clknet_leaf_65_clk _0447_ VGND VGND VPWR VPWR rf.registers\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6499_ net13 net12 net11 VGND VGND VPWR VPWR _3153_ sky130_fd_sc_hd__or3_4
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7092__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7485__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5605__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8238_ net274 _3450_ _4060_ VGND VGND VPWR VPWR _4094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4394__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8169_ _4057_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7788__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4697__S1 _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6870__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_41_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7206__S _3539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4385__S0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7779__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5239__C1 _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6451__A1 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5870_ _2246_ _2616_ VGND VGND VPWR VPWR _2617_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4821_ rf.registers\[20\]\[16\] rf.registers\[21\]\[16\] rf.registers\[22\]\[16\]
+ rf.registers\[23\]\[16\] _1291_ _1194_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7951__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7540_ _3724_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
X_4752_ rf.registers\[0\]\[15\] rf.registers\[1\]\[15\] rf.registers\[2\]\[15\] rf.registers\[3\]\[15\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_78_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7471_ _3067_ net899 _3686_ VGND VGND VPWR VPWR _3688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4683_ _1189_ _1438_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6422_ net41 VGND VGND VPWR VPWR _3103_ sky130_fd_sc_hd__buf_2
X_9210_ clknet_leaf_35_clk _0370_ VGND VGND VPWR VPWR rf.registers\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8500__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9141_ clknet_leaf_38_clk _0301_ VGND VGND VPWR VPWR rf.registers\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6353_ _3055_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5304_ _2058_ _2059_ _1685_ VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9072_ clknet_leaf_3_clk _0232_ VGND VGND VPWR VPWR rf.registers\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6284_ net407 _3002_ _3007_ VGND VGND VPWR VPWR _3008_ sky130_fd_sc_hd__mux2_1
X_8023_ _3145_ net1022 _3974_ VGND VGND VPWR VPWR _3980_ sky130_fd_sc_hd__mux2_1
X_5235_ rf.registers\[4\]\[26\] rf.registers\[5\]\[26\] rf.registers\[6\]\[26\] rf.registers\[7\]\[26\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__mux4_1
XANTENNA__4376__S0 _1065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5166_ _1766_ _1921_ _1672_ VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__o21ai_1
X_5097_ _1700_ _1852_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5160__A _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6442__A1 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4679__S1 _1184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8925_ clknet_leaf_15_clk _0085_ VGND VGND VPWR VPWR rf.registers\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6690__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8856_ clknet_leaf_27_clk _0016_ VGND VGND VPWR VPWR rf.registers\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7807_ _3865_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__clkbuf_1
X_5999_ _2585_ _2738_ _2333_ VGND VGND VPWR VPWR _2739_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7942__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8787_ clknet_leaf_33_clk _0971_ VGND VGND VPWR VPWR rf.registers\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7738_ _3062_ net1152 _3819_ VGND VGND VPWR VPWR _3829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4851__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7669_ _3792_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9408_ clknet_leaf_60_clk _0568_ VGND VGND VPWR VPWR rf.registers\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5181__A1 _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9339_ clknet_leaf_34_clk _0499_ VGND VGND VPWR VPWR rf.registers\[21\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7458__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7026__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6865__S _3340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6681__A1 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8186__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5095__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4414__A _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4842__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8320__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold409 rf.registers\[17\]\[27\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4358__S0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5020_ _1774_ _1775_ _1726_ VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_2_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7621__A0 _3081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6971_ net1045 _3009_ _3398_ VGND VGND VPWR VPWR _3406_ sky130_fd_sc_hd__mux2_1
X_8710_ clknet_leaf_5_clk _0894_ VGND VGND VPWR VPWR rf.registers\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5922_ _2193_ _2640_ _2641_ VGND VGND VPWR VPWR _2666_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8641_ clknet_leaf_56_clk _0825_ VGND VGND VPWR VPWR rf.registers\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5853_ _2539_ _2559_ _2560_ VGND VGND VPWR VPWR _2601_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_152_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7924__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4804_ rf.registers\[28\]\[11\] rf.registers\[29\]\[11\] rf.registers\[30\]\[11\]
+ rf.registers\[31\]\[11\] _1042_ _1044_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__mux4_2
XANTENNA__4738__A1 _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5784_ _2534_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_1
X_8572_ clknet_leaf_16_clk _0756_ VGND VGND VPWR VPWR rf.registers\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4833__S1 _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7523_ _3715_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
X_4735_ rf.registers\[12\]\[14\] rf.registers\[13\]\[14\] rf.registers\[14\]\[14\]
+ rf.registers\[15\]\[14\] net1156 _1279_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7454_ _3050_ net171 _3675_ VGND VGND VPWR VPWR _3679_ sky130_fd_sc_hd__mux2_1
XANTENNA__8230__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4666_ rf.registers\[8\]\[23\] rf.registers\[9\]\[23\] rf.registers\[10\]\[23\] rf.registers\[11\]\[23\]
+ net1164 _1268_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6405_ net10 net9 net46 VGND VGND VPWR VPWR _3091_ sky130_fd_sc_hd__nand3b_4
XANTENNA__4597__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7385_ _3642_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
Xhold910 rf.registers\[21\]\[20\] VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold921 rf.registers\[17\]\[9\] VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__dlygate4sd3_1
X_4597_ rf.registers\[20\]\[25\] rf.registers\[21\]\[25\] rf.registers\[22\]\[25\]
+ rf.registers\[23\]\[25\] _1351_ _1352_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__mux4_1
Xhold932 rf.registers\[13\]\[14\] VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold943 rf.registers\[14\]\[22\] VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__dlygate4sd3_1
X_9124_ clknet_leaf_47_clk _0284_ VGND VGND VPWR VPWR rf.registers\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6336_ _3022_ VGND VGND VPWR VPWR _3044_ sky130_fd_sc_hd__clkbuf_8
Xhold954 rf.registers\[12\]\[26\] VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 rf.registers\[4\]\[8\] VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 rf.registers\[30\]\[22\] VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 rf.registers\[2\]\[15\] VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__dlygate4sd3_1
X_9055_ clknet_leaf_74_clk _0215_ VGND VGND VPWR VPWR rf.registers\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold998 rf.registers\[14\]\[31\] VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__dlygate4sd3_1
X_6267_ net92 _2981_ _2741_ VGND VGND VPWR VPWR _2992_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6663__A1 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8006_ _3128_ net600 _3963_ VGND VGND VPWR VPWR _3971_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5218_ rf.registers\[4\]\[27\] rf.registers\[5\]\[27\] rf.registers\[6\]\[27\] rf.registers\[7\]\[27\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__mux4_1
X_6198_ _2530_ _2792_ _2922_ _2926_ VGND VGND VPWR VPWR _2927_ sky130_fd_sc_hd__o211a_1
X_5149_ _1842_ _1904_ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8405__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8908_ clknet_leaf_45_clk _0068_ VGND VGND VPWR VPWR rf.registers\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8168__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8839_ clknet_leaf_1_clk _1023_ VGND VGND VPWR VPWR rf.registers\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7915__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4824__S1 _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4674__A1_N _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4588__S0 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6595__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6654__A1 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4760__S0 _1026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4843__S _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5068__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5917__B1 _2175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8050__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4520_ _1254_ _1275_ _1171_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold206 rf.registers\[10\]\[9\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _1191_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__buf_12
XFILLER_0_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold217 rf.registers\[6\]\[20\] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4579__S0 _1267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold228 rf.registers\[5\]\[3\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold239 rf.registers\[3\]\[12\] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
X_7170_ net162 _3474_ _3517_ VGND VGND VPWR VPWR _3527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4382_ _1136_ _1137_ _1047_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6121_ _1731_ _2853_ VGND VGND VPWR VPWR _2854_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6052_ _2421_ _2788_ VGND VGND VPWR VPWR _2789_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5003_ rf.registers\[20\]\[21\] rf.registers\[21\]\[21\] rf.registers\[22\]\[21\]
+ rf.registers\[23\]\[21\] _1676_ _1681_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4751__S0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8398__A1 _3474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4753__S _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6954_ net311 _3132_ _3387_ VGND VGND VPWR VPWR _3397_ sky130_fd_sc_hd__mux2_1
XANTENNA__5081__B1 _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5905_ _2609_ _2649_ _1803_ VGND VGND VPWR VPWR _2650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6885_ _3360_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8624_ clknet_leaf_4_clk _0808_ VGND VGND VPWR VPWR rf.registers\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_5836_ _2579_ _2583_ _2252_ VGND VGND VPWR VPWR _2584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4806__S1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5767_ _2516_ _2517_ VGND VGND VPWR VPWR _2518_ sky130_fd_sc_hd__nor2_1
X_8555_ _4261_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4989__A _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7506_ _3706_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
X_4718_ _1472_ _1473_ _1287_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8322__A1 _3466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5698_ _2449_ _2451_ VGND VGND VPWR VPWR _2452_ sky130_fd_sc_hd__nand2_1
X_8486_ _4225_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__clkbuf_1
X_4649_ _1403_ _1404_ _1107_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__mux2_1
X_7437_ _3033_ net550 _3664_ VGND VGND VPWR VPWR _3670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold740 rf.registers\[11\]\[19\] VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__dlygate4sd3_1
X_7368_ _3633_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
Xhold751 rf.registers\[31\]\[7\] VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold762 rf.registers\[24\]\[28\] VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 rf.registers\[4\]\[17\] VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd3_1
X_9107_ clknet_leaf_34_clk _0267_ VGND VGND VPWR VPWR rf.registers\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6319_ _3032_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8196__A _4060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold784 rf.registers\[3\]\[31\] VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd3_1
X_7299_ _3596_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6709__A _3266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4990__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold795 rf.registers\[31\]\[21\] VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7304__S _3591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5613__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9038_ clknet_leaf_43_clk _0198_ VGND VGND VPWR VPWR rf.registers\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8135__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5298__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6444__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__8010__A0 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4899__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5494__S _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5470__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4981__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7214__S _3516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4638__B1 _1037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6354__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5063__B1 _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6670_ _3246_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8552__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5621_ _2335_ _2337_ _2340_ _2375_ _2333_ VGND VGND VPWR VPWR _2376_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_14_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5366__B2 _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5552_ rf.registers\[20\]\[5\] rf.registers\[21\]\[5\] rf.registers\[22\]\[5\] rf.registers\[23\]\[5\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2308_ sky130_fd_sc_hd__mux4_1
XANTENNA__5461__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8340_ _4148_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4503_ _1036_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8271_ _3120_ net276 _4108_ VGND VGND VPWR VPWR _4112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5483_ rf.registers\[8\]\[9\] rf.registers\[9\]\[9\] rf.registers\[10\]\[9\] rf.registers\[11\]\[9\]
+ _1782_ _1692_ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7222_ _3019_ net567 _3555_ VGND VGND VPWR VPWR _3556_ sky130_fd_sc_hd__mux2_1
X_4434_ _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4877__B1 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7153_ _3518_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_4365_ rf.registers\[8\]\[2\] rf.registers\[9\]\[2\] rf.registers\[10\]\[2\] rf.registers\[11\]\[2\]
+ net101 _1066_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7124__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6104_ _1754_ _2837_ VGND VGND VPWR VPWR _2838_ sky130_fd_sc_hd__nand2_1
X_7084_ _3473_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
X_4296_ net93 VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__buf_12
XANTENNA__5826__C1 _2373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6035_ _1858_ _2762_ _2772_ VGND VGND VPWR VPWR _2773_ sky130_fd_sc_hd__a21o_1
XANTENNA__6963__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer10 net91 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer32 _1528_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer43 net124 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer54 _2885_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlymetal6s2s_1
X_7986_ _3960_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__clkbuf_1
X_6937_ _3388_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_36_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7794__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4801__B1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6868_ net200 _3113_ _3351_ VGND VGND VPWR VPWR _3352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8607_ clknet_leaf_73_clk _0791_ VGND VGND VPWR VPWR rf.registers\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5819_ _2458_ _2567_ _1126_ VGND VGND VPWR VPWR _2568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9587_ clknet_leaf_32_clk _0747_ VGND VGND VPWR VPWR rf.registers\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6799_ _3303_ VGND VGND VPWR VPWR _3315_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__7095__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8538_ _4252_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8469_ net355 net15 _4216_ VGND VGND VPWR VPWR _4217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6857__A1 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold570 rf.registers\[2\]\[1\] VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 rf.registers\[24\]\[15\] VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7034__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold592 rf.registers\[5\]\[0\] VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5343__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6174__A _1996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5045__B1 _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5443__S1 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4422__A _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4954__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_50_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7879__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6783__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7840_ _3883_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6233__C1 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7771_ net451 _3460_ _3844_ VGND VGND VPWR VPWR _3847_ sky130_fd_sc_hd__mux2_1
XANTENNA__5131__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4983_ _1738_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__clkbuf_8
X_9510_ clknet_leaf_66_clk _0670_ VGND VGND VPWR VPWR rf.registers\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6722_ _3035_ net729 _3267_ VGND VGND VPWR VPWR _3274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8525__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9441_ clknet_leaf_61_clk _0601_ VGND VGND VPWR VPWR rf.registers\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6653_ _3237_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5434__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4332__A _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5604_ _2357_ _2358_ VGND VGND VPWR VPWR _2359_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9372_ clknet_leaf_17_clk _0532_ VGND VGND VPWR VPWR rf.registers\[20\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6584_ _3033_ net1107 _3195_ VGND VGND VPWR VPWR _3201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8323_ _4139_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5535_ rf.registers\[16\]\[4\] rf.registers\[17\]\[4\] rf.registers\[18\]\[4\] rf.registers\[19\]\[4\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6839__A1 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5198__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8254_ _3103_ net437 _4097_ VGND VGND VPWR VPWR _4103_ sky130_fd_sc_hd__mux2_1
X_5466_ rf.registers\[12\]\[8\] rf.registers\[13\]\[8\] rf.registers\[14\]\[8\] rf.registers\[15\]\[8\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4417_ net1156 VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__buf_12
X_7205_ _3545_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
X_8185_ _4066_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__clkbuf_1
X_5397_ _1684_ _2152_ VGND VGND VPWR VPWR _2153_ sky130_fd_sc_hd__or2_1
XANTENNA__6259__A _1923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5163__A _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7136_ net484 _3508_ _3498_ VGND VGND VPWR VPWR _3509_ sky130_fd_sc_hd__mux2_1
X_4348_ _1041_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__buf_12
X_7067_ net39 VGND VGND VPWR VPWR _3462_ sky130_fd_sc_hd__buf_2
X_4279_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__buf_4
X_6018_ _2527_ _2756_ _2426_ VGND VGND VPWR VPWR _2757_ sky130_fd_sc_hd__mux2_1
XANTENNA__5370__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4507__A _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7969_ _3021_ _3552_ VGND VGND VPWR VPWR _3951_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_120_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8413__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8516__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5425__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6868__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5189__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7699__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7007__A1 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4417__A net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5416__S1 _1721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer1 _1125_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_70_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5320_ rf.registers\[4\]\[2\] rf.registers\[5\]\[2\] rf.registers\[6\]\[2\] rf.registers\[7\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2076_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5251_ rf.registers\[8\]\[25\] rf.registers\[9\]\[25\] rf.registers\[10\]\[25\] rf.registers\[11\]\[25\]
+ _1895_ _1897_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__mux4_1
XANTENNA__4927__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5182_ rf.registers\[8\]\[29\] rf.registers\[9\]\[29\] rf.registers\[10\]\[29\] rf.registers\[11\]\[29\]
+ _1767_ _1768_ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8941_ clknet_leaf_44_clk _0101_ VGND VGND VPWR VPWR rf.registers\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5352__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8872_ clknet_leaf_47_clk _0032_ VGND VGND VPWR VPWR rf.registers\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_7823_ net854 _3444_ _3866_ VGND VGND VPWR VPWR _3874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7754_ _3837_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4966_ _1721_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__buf_4
X_6705_ _3264_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7685_ net188 _3442_ _3794_ VGND VGND VPWR VPWR _3801_ sky130_fd_sc_hd__mux2_1
X_4897_ _1651_ _1652_ net3 VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5407__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9424_ clknet_leaf_11_clk _0584_ VGND VGND VPWR VPWR rf.registers\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6636_ _3085_ net1127 _3194_ VGND VGND VPWR VPWR _3228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9355_ clknet_leaf_4_clk _0515_ VGND VGND VPWR VPWR rf.registers\[20\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6688__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6567_ _3190_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8306_ _3015_ net389 _4096_ VGND VGND VPWR VPWR _4130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5518_ rf.registers\[28\]\[7\] rf.registers\[29\]\[7\] rf.registers\[30\]\[7\] rf.registers\[31\]\[7\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2274_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9286_ clknet_leaf_72_clk _0446_ VGND VGND VPWR VPWR rf.registers\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6498_ _3152_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__clkbuf_1
X_8237_ _4093_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__clkbuf_1
X_5449_ _1699_ _2204_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__nand2_1
X_8168_ net547 _3448_ _4047_ VGND VGND VPWR VPWR _4057_ sky130_fd_sc_hd__mux2_1
XANTENNA__4394__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7119_ net26 VGND VGND VPWR VPWR _3497_ sky130_fd_sc_hd__clkbuf_4
X_8099_ _4020_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8143__S _4036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5420__B1 _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_rebuffer51_A _1277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8379__A _4168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4385__S1 _1090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8318__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7222__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5531__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6739__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5677__S _2363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4820_ rf.registers\[16\]\[16\] rf.registers\[17\]\[16\] rf.registers\[18\]\[16\]
+ rf.registers\[19\]\[16\] _1291_ _1194_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4751_ rf.registers\[4\]\[15\] rf.registers\[5\]\[15\] rf.registers\[6\]\[15\] rf.registers\[7\]\[15\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7470_ _3687_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
X_4682_ rf.registers\[8\]\[22\] rf.registers\[9\]\[22\] rf.registers\[10\]\[22\] rf.registers\[11\]\[22\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__mux4_1
XFILLER_0_141_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6421_ _3102_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5714__A1 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7193__A _3516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9140_ clknet_leaf_42_clk _0300_ VGND VGND VPWR VPWR rf.registers\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6352_ _3054_ net950 _3044_ VGND VGND VPWR VPWR _3055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5303_ rf.registers\[0\]\[3\] rf.registers\[1\]\[3\] rf.registers\[2\]\[3\] rf.registers\[3\]\[3\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__mux4_1
X_9071_ clknet_leaf_8_clk _0231_ VGND VGND VPWR VPWR rf.registers\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6283_ _3006_ VGND VGND VPWR VPWR _3007_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8022_ _3979_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__clkbuf_1
X_5234_ _1988_ _1989_ _1901_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__mux2_1
XANTENNA__4376__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8228__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5165_ _1917_ _1920_ _1901_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5096_ _1850_ _1851_ _1713_ VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__mux2_1
XANTENNA__6971__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8924_ clknet_leaf_18_clk _0084_ VGND VGND VPWR VPWR rf.registers\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8855_ clknet_leaf_24_clk _0015_ VGND VGND VPWR VPWR rf.registers\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7806_ net360 _3495_ _3855_ VGND VGND VPWR VPWR _3865_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8786_ clknet_leaf_25_clk _0970_ VGND VGND VPWR VPWR rf.registers\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5998_ _1127_ _2737_ VGND VGND VPWR VPWR _2738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7737_ _3828_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__clkbuf_1
X_4949_ _1704_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__buf_4
XFILLER_0_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_rebuffer1_A _1125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7668_ net339 _3493_ _3783_ VGND VGND VPWR VPWR _3792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9407_ clknet_leaf_71_clk _0567_ VGND VGND VPWR VPWR rf.registers\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6619_ _3219_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7599_ _3755_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9338_ clknet_leaf_35_clk _0498_ VGND VGND VPWR VPWR rf.registers\[21\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9269_ clknet_leaf_31_clk _0429_ VGND VGND VPWR VPWR rf.registers\[23\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6130__A1 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5564__S0 _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6447__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7042__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5316__S0 _1701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7977__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6197__A1 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4358__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5555__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4576__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8048__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6357__A net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5261__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7887__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6791__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6970_ _3405_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5921_ _2598_ _2617_ _2664_ VGND VGND VPWR VPWR _2665_ sky130_fd_sc_hd__nand3_2
XFILLER_0_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8640_ clknet_leaf_68_clk _0824_ VGND VGND VPWR VPWR rf.registers\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4605__A _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5852_ _2511_ _2512_ _2518_ _2542_ _2599_ VGND VGND VPWR VPWR _2600_ sky130_fd_sc_hd__a311o_1
XANTENNA__5200__S _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4803_ rf.registers\[24\]\[11\] rf.registers\[25\]\[11\] rf.registers\[26\]\[11\]
+ rf.registers\[27\]\[11\] _1072_ _1073_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__mux4_2
X_8571_ clknet_leaf_21_clk _0755_ VGND VGND VPWR VPWR rf.registers\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5783_ _2521_ _2529_ _2533_ VGND VGND VPWR VPWR _2534_ sky130_fd_sc_hd__or3_1
XFILLER_0_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7522_ _3050_ net372 _3711_ VGND VGND VPWR VPWR _3715_ sky130_fd_sc_hd__mux2_1
X_4734_ rf.registers\[8\]\[14\] rf.registers\[9\]\[14\] rf.registers\[10\]\[14\] rf.registers\[11\]\[14\]
+ net1161 _1279_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__mux4_1
XANTENNA__6820__A _3303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7453_ _3678_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _1417_ _1418_ _1419_ _1420_ _1190_ _1205_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7127__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6404_ net12 net11 net13 VGND VGND VPWR VPWR _3090_ sky130_fd_sc_hd__or3b_4
Xhold900 rf.registers\[21\]\[5\] VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold911 rf.registers\[6\]\[13\] VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__dlygate4sd3_1
X_7384_ _3048_ net1018 _3639_ VGND VGND VPWR VPWR _3642_ sky130_fd_sc_hd__mux2_1
XANTENNA__4597__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold922 rf.registers\[13\]\[4\] VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4596_ _1325_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__clkbuf_4
X_9123_ clknet_leaf_68_clk _0283_ VGND VGND VPWR VPWR rf.registers\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold933 rf.registers\[26\]\[27\] VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold944 rf.registers\[25\]\[6\] VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__dlygate4sd3_1
X_6335_ net15 VGND VGND VPWR VPWR _3043_ sky130_fd_sc_hd__clkbuf_2
Xhold955 rf.registers\[20\]\[2\] VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 rf.registers\[8\]\[2\] VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7651__A _3771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold977 rf.registers\[8\]\[27\] VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__dlygate4sd3_1
X_9054_ clknet_leaf_74_clk _0214_ VGND VGND VPWR VPWR rf.registers\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold988 rf.registers\[20\]\[14\] VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5546__S0 _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold999 rf.registers\[3\]\[10\] VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__dlygate4sd3_1
X_6266_ _2952_ _2986_ _2987_ _2984_ VGND VGND VPWR VPWR _2991_ sky130_fd_sc_hd__a31o_1
X_8005_ _3970_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4486__S _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8979__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5217_ _1773_ _1972_ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_110_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6197_ _2337_ _2925_ _1086_ VGND VGND VPWR VPWR _2926_ sky130_fd_sc_hd__o21a_1
X_5148_ _1777_ _1890_ _1894_ _1903_ VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_86_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5079_ rf.registers\[0\]\[19\] rf.registers\[1\]\[19\] rf.registers\[2\]\[19\] rf.registers\[3\]\[19\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__mux4_1
X_8907_ clknet_leaf_4_clk _0067_ VGND VGND VPWR VPWR rf.registers\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7098__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8838_ clknet_leaf_1_clk _1022_ VGND VGND VPWR VPWR rf.registers\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8769_ clknet_leaf_56_clk _0953_ VGND VGND VPWR VPWR rf.registers\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6730__A _3266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7679__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5346__A _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4588__S1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5065__B _1820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6876__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5537__S0 _2050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4396__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6177__A _2626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4760__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4425__A _1042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5020__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4276__S0 _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4450_ _1199_ _1204_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__a21o_1
Xhold207 rf.registers\[6\]\[5\] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4579__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold218 rf.registers\[11\]\[3\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold229 rf.registers\[4\]\[19\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4353__B1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4381_ rf.registers\[12\]\[1\] rf.registers\[13\]\[1\] rf.registers\[14\]\[1\] rf.registers\[15\]\[1\]
+ net117 _1053_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6120_ _1430_ _2852_ VGND VGND VPWR VPWR _2853_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6051_ _2784_ _2787_ VGND VGND VPWR VPWR _2788_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5002_ _1639_ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4751__S1 _1195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8506__S _4227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6953_ _3396_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5081__A1 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5904_ _2352_ _2350_ VGND VGND VPWR VPWR _2649_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6884_ net489 _3130_ _3351_ VGND VGND VPWR VPWR _3360_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_81_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8623_ clknet_leaf_10_clk _0807_ VGND VGND VPWR VPWR rf.registers\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_5835_ _2547_ _2582_ _2363_ VGND VGND VPWR VPWR _2583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8554_ net903 net24 _4255_ VGND VGND VPWR VPWR _4261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5766_ _2323_ _2515_ VGND VGND VPWR VPWR _2517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7505_ _3033_ net671 _3700_ VGND VGND VPWR VPWR _3706_ sky130_fd_sc_hd__mux2_1
X_4717_ rf.registers\[12\]\[13\] rf.registers\[13\]\[13\] rf.registers\[14\]\[13\]
+ rf.registers\[15\]\[13\] _1291_ _1194_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__mux4_1
X_8485_ net847 net23 _4216_ VGND VGND VPWR VPWR _4225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5697_ _2450_ _2414_ _2413_ VGND VGND VPWR VPWR _2451_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_115_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7436_ _3669_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_1
X_4648_ rf.registers\[24\]\[7\] rf.registers\[25\]\[7\] rf.registers\[26\]\[7\] rf.registers\[27\]\[7\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1 _1181_ VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_96_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6696__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold730 rf.registers\[29\]\[23\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
X_7367_ _3031_ net738 _3628_ VGND VGND VPWR VPWR _3633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold741 rf.registers\[30\]\[17\] VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd3_1
X_4579_ rf.registers\[24\]\[30\] rf.registers\[25\]\[30\] rf.registers\[26\]\[30\]
+ rf.registers\[27\]\[30\] _1267_ _1268_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold752 rf.registers\[24\]\[26\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd3_1
X_9106_ clknet_leaf_39_clk _0266_ VGND VGND VPWR VPWR rf.registers\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8086__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold763 rf.registers\[24\]\[21\] VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ _3031_ net510 _3023_ VGND VGND VPWR VPWR _3032_ sky130_fd_sc_hd__mux2_1
Xhold774 rf.registers\[26\]\[19\] VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5519__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold785 rf.registers\[30\]\[15\] VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd3_1
X_7298_ _3031_ net530 _3591_ VGND VGND VPWR VPWR _3596_ sky130_fd_sc_hd__mux2_1
Xhold796 rf.registers\[18\]\[30\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4990__S1 _1723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9037_ clknet_leaf_50_clk _0197_ VGND VGND VPWR VPWR rf.registers\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6249_ _1148_ _1925_ VGND VGND VPWR VPWR _2975_ sky130_fd_sc_hd__nand2_1
XANTENNA__5844__B1 _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8077__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4981__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5015__S _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4638__A1 _1036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8326__S _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7230__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold90 rf.registers\[18\]\[9\] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5063__A1 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8061__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5620_ _2105_ _2356_ _2374_ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__o21ai_1
XANTENNA__6370__A net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ _1799_ _2306_ VGND VGND VPWR VPWR _2307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4502_ rf.registers\[16\]\[21\] rf.registers\[17\]\[21\] rf.registers\[18\]\[21\]
+ rf.registers\[19\]\[21\] _1220_ _1222_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__mux4_2
X_8270_ _4111_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__clkbuf_1
X_5482_ rf.registers\[12\]\[9\] rf.registers\[13\]\[9\] rf.registers\[14\]\[9\] rf.registers\[15\]\[9\]
+ _1782_ _1680_ VGND VGND VPWR VPWR _2238_ sky130_fd_sc_hd__mux4_1
XANTENNA__4326__B1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7221_ _3554_ VGND VGND VPWR VPWR _3555_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4433_ _1048_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__buf_4
XANTENNA__4877__A1 _1254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4421__S0 _1173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7405__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7152_ net346 _3454_ _3517_ VGND VGND VPWR VPWR _3518_ sky130_fd_sc_hd__mux2_1
X_4364_ _1047_ _1119_ _1050_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6103_ _1446_ _2836_ VGND VGND VPWR VPWR _2837_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7815__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4295_ _1048_ _1049_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__o21a_1
X_7083_ net220 _3472_ _3456_ VGND VGND VPWR VPWR _3473_ sky130_fd_sc_hd__mux2_1
X_6034_ _1874_ _2743_ _2762_ _1858_ VGND VGND VPWR VPWR _2772_ sky130_fd_sc_hd__o22a_1
XANTENNA__8236__S _4083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6545__A _3156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7140__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer11 _1238_ VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer22 _1256_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer33 net114 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer44 _2657_ VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__dlymetal6s2s_1
X_7985_ _3107_ net328 _3952_ VGND VGND VPWR VPWR _3960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4488__S0 _1207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6936_ net609 _3113_ _3387_ VGND VGND VPWR VPWR _3388_ sky130_fd_sc_hd__mux2_1
XANTENNA__4801__A1 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6867_ _3339_ VGND VGND VPWR VPWR _3351_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8606_ clknet_leaf_73_clk _0790_ VGND VGND VPWR VPWR rf.registers\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5818_ _2525_ _2566_ _1146_ VGND VGND VPWR VPWR _2567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7751__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9586_ clknet_leaf_27_clk _0746_ VGND VGND VPWR VPWR rf.registers\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6798_ _3314_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8537_ net221 net16 _4244_ VGND VGND VPWR VPWR _4252_ sky130_fd_sc_hd__mux2_1
X_5749_ _1126_ VGND VGND VPWR VPWR _2501_ sky130_fd_sc_hd__clkbuf_4
X_8468_ _4204_ VGND VGND VPWR VPWR _4216_ sky130_fd_sc_hd__buf_4
X_7419_ _3083_ net832 _3650_ VGND VGND VPWR VPWR _3660_ sky130_fd_sc_hd__mux2_1
XANTENNA__4939__S _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8399_ _4179_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7315__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5624__A _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold560 rf.registers\[6\]\[14\] VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold571 rf.registers\[14\]\[24\] VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 rf.registers\[18\]\[15\] VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 rf.registers\[12\]\[24\] VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7806__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7985__S _3952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6793__A1 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4651__S0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4849__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4403__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4954__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output72_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput80 net80 VGND VGND VPWR VPWR alu_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_128_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5808__B1 _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8056__S _3989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8222__A1 _3502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7895__S _3902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7770_ _3846_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__clkbuf_1
X_4982_ _1684_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__7981__A0 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5131__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6721_ _3273_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9440_ clknet_leaf_69_clk _0600_ VGND VGND VPWR VPWR rf.registers\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6652_ rf.registers\[8\]\[5\] _3103_ _3231_ VGND VGND VPWR VPWR _3237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5603_ _1839_ _2230_ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9371_ clknet_leaf_34_clk _0531_ VGND VGND VPWR VPWR rf.registers\[20\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6583_ _3200_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8322_ net930 _3466_ _4133_ VGND VGND VPWR VPWR _4139_ sky130_fd_sc_hd__mux2_1
X_5534_ rf.registers\[20\]\[4\] rf.registers\[21\]\[4\] rf.registers\[22\]\[4\] rf.registers\[23\]\[4\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2290_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8253_ _4102_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4759__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5465_ rf.registers\[8\]\[8\] rf.registers\[9\]\[8\] rf.registers\[10\]\[8\] rf.registers\[11\]\[8\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _2221_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_76_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5198__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7204_ net507 _3508_ _3539_ VGND VGND VPWR VPWR _3545_ sky130_fd_sc_hd__mux2_1
X_4416_ _1072_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__buf_12
XFILLER_0_111_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8184_ net319 _3464_ _4061_ VGND VGND VPWR VPWR _4066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5396_ rf.registers\[4\]\[13\] rf.registers\[5\]\[13\] rf.registers\[6\]\[13\] rf.registers\[7\]\[13\]
+ _1702_ _1678_ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7135_ net31 VGND VGND VPWR VPWR _3508_ sky130_fd_sc_hd__buf_2
X_4347_ rf.registers\[4\]\[3\] rf.registers\[5\]\[3\] rf.registers\[6\]\[3\] rf.registers\[7\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__mux4_1
X_7066_ _3461_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
X_4278_ net6 VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__inv_2
X_6017_ _2565_ _2609_ _1148_ VGND VGND VPWR VPWR _2756_ sky130_fd_sc_hd__mux2_1
XANTENNA__5370__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8213__A1 _3493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ _3950_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919_ net871 _3097_ _3376_ VGND VGND VPWR VPWR _3379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7899_ _3017_ net915 _3879_ VGND VGND VPWR VPWR _3914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4523__A _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6527__A1 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9569_ clknet_leaf_67_clk _0729_ VGND VGND VPWR VPWR rf.registers\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4633__S0 _1219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7834__A _3879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5189__S1 _1884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7045__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold390 rf.registers\[10\]\[15\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6884__S _3351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8452__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6215__B1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6518__A1 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4433__A _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7191__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5963__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4624__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_20_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer2 net83 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5741__A2 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5250_ _2002_ _2005_ _1700_ VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__mux2_1
XANTENNA__4927__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5181_ _1745_ _1936_ _1697_ VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_71_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8940_ clknet_leaf_45_clk _0100_ VGND VGND VPWR VPWR rf.registers\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6095__A _1779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5352__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8871_ clknet_leaf_65_clk _0031_ VGND VGND VPWR VPWR rf.registers\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7822_ _3873_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8514__S _3007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7753_ _3077_ net756 _3830_ VGND VGND VPWR VPWR _3837_ sky130_fd_sc_hd__mux2_1
X_4965_ _1678_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6704_ net318 _3015_ _3230_ VGND VGND VPWR VPWR _3264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7684_ _3800_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__clkbuf_1
X_4896_ rf.registers\[12\]\[0\] rf.registers\[13\]\[0\] rf.registers\[14\]\[0\] rf.registers\[15\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5980__A2 _2530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9423_ clknet_leaf_28_clk _0583_ VGND VGND VPWR VPWR rf.registers\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6635_ _3227_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6969__S _3398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9354_ clknet_leaf_63_clk _0514_ VGND VGND VPWR VPWR rf.registers\[20\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6566_ net566 _3015_ _3156_ VGND VGND VPWR VPWR _3190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8305_ _4129_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__clkbuf_1
X_5517_ rf.registers\[24\]\[7\] rf.registers\[25\]\[7\] rf.registers\[26\]\[7\] rf.registers\[27\]\[7\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2273_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4489__S _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9285_ clknet_leaf_57_clk _0445_ VGND VGND VPWR VPWR rf.registers\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6497_ net159 _3017_ _3092_ VGND VGND VPWR VPWR _3152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8236_ net525 _3448_ _4083_ VGND VGND VPWR VPWR _4093_ sky130_fd_sc_hd__mux2_1
X_5448_ _2202_ _2203_ _1711_ VGND VGND VPWR VPWR _2204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8167_ _4056_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__clkbuf_1
X_5379_ _1699_ _2134_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__nand2_1
XANTENNA__8434__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7118_ _3496_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_8098_ net1147 _3446_ _4011_ VGND VGND VPWR VPWR _4020_ sky130_fd_sc_hd__mux2_1
X_7049_ _3449_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6996__A1 _3105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8424__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5349__A _2104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4854__S0 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7173__A1 _3476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5031__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7503__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5239__A1 _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5531__B _2286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4428__A _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__S0 _1822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4750_ _1214_ _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6789__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7164__A1 _3468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4681_ _1433_ _1436_ _1187_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6420_ net250 _3101_ _3093_ VGND VGND VPWR VPWR _3102_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6351_ net20 VGND VGND VPWR VPWR _3054_ sky130_fd_sc_hd__buf_2
XFILLER_0_52_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5302_ rf.registers\[4\]\[3\] rf.registers\[5\]\[3\] rf.registers\[6\]\[3\] rf.registers\[7\]\[3\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_73_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9070_ clknet_leaf_41_clk _0230_ VGND VGND VPWR VPWR rf.registers\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6282_ _3003_ _3005_ VGND VGND VPWR VPWR _3006_ sky130_fd_sc_hd__nor2_4
XFILLER_0_122_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8021_ _3143_ net651 _3974_ VGND VGND VPWR VPWR _3979_ sky130_fd_sc_hd__mux2_1
X_5233_ rf.registers\[8\]\[26\] rf.registers\[9\]\[26\] rf.registers\[10\]\[26\] rf.registers\[11\]\[26\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7413__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8608__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5164_ rf.registers\[0\]\[30\] rf.registers\[1\]\[30\] rf.registers\[2\]\[30\] rf.registers\[3\]\[30\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__mux4_1
XANTENNA__4338__A _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5095_ rf.registers\[12\]\[17\] rf.registers\[13\]\[17\] rf.registers\[14\]\[17\]
+ rf.registers\[15\]\[17\] _1720_ _1723_ VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__mux4_1
X_8923_ clknet_leaf_22_clk _0083_ VGND VGND VPWR VPWR rf.registers\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8244__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8854_ clknet_leaf_24_clk _0014_ VGND VGND VPWR VPWR rf.registers\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7805_ _3864_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__clkbuf_1
X_8785_ clknet_leaf_44_clk _0969_ VGND VGND VPWR VPWR rf.registers\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _1060_ _1085_ VGND VGND VPWR VPWR _2737_ sky130_fd_sc_hd__nor2b_2
XANTENNA__4836__S0 _1287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5169__A _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7736_ _3060_ net1039 _3819_ VGND VGND VPWR VPWR _3828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4948_ _1703_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7667_ _3791_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
X_4879_ _1602_ _1618_ _1634_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5166__B1 _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9406_ clknet_leaf_72_clk _0566_ VGND VGND VPWR VPWR rf.registers\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6618_ _3067_ net765 _3217_ VGND VGND VPWR VPWR _3219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7598_ _3058_ net897 _3747_ VGND VGND VPWR VPWR _3755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6549_ _3181_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__clkbuf_1
X_9337_ clknet_leaf_20_clk _0497_ VGND VGND VPWR VPWR rf.registers\[21\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9268_ clknet_leaf_42_clk _0428_ VGND VGND VPWR VPWR rf.registers\[23\]\[22\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5013__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8219_ _4084_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8419__S _4180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9199_ clknet_leaf_9_clk _0359_ VGND VGND VPWR VPWR rf.registers\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5564__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7323__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_144_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5316__S1 _1677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8154__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4827__S0 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5252__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5004__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5555__S1 _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5880__B2 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5632__A1 _1168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5920_ _2633_ _2642_ _2643_ VGND VGND VPWR VPWR _2664_ sky130_fd_sc_hd__and3_1
XANTENNA__6373__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5851_ _2562_ _2560_ _2559_ VGND VGND VPWR VPWR _2599_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4818__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4802_ _1024_ _1549_ _1553_ _1557_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__a2bb2o_4
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8570_ clknet_leaf_18_clk _0754_ VGND VGND VPWR VPWR rf.registers\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5782_ _2530_ _2531_ _2532_ _2373_ VGND VGND VPWR VPWR _2533_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7521_ _3714_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4733_ _1287_ _1488_ _1078_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6312__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7452_ _3048_ net868 _3675_ VGND VGND VPWR VPWR _3678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4664_ rf.registers\[20\]\[23\] rf.registers\[21\]\[23\] rf.registers\[22\]\[23\]
+ rf.registers\[23\]\[23\] _1351_ _1352_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6403_ net14 VGND VGND VPWR VPWR _3089_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7383_ _3641_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
Xhold901 rf.registers\[1\]\[7\] VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__dlygate4sd3_1
X_4595_ _1324_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__buf_8
Xhold912 rf.registers\[16\]\[10\] VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9122_ clknet_leaf_58_clk _0282_ VGND VGND VPWR VPWR rf.registers\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold923 rf.registers\[23\]\[1\] VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6334_ _3042_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__clkbuf_1
Xhold934 rf.registers\[23\]\[24\] VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 rf.registers\[15\]\[23\] VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 rf.registers\[22\]\[6\] VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 rf.registers\[24\]\[24\] VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold978 rf.registers\[27\]\[9\] VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__dlygate4sd3_1
X_9053_ clknet_leaf_15_clk _0213_ VGND VGND VPWR VPWR rf.registers\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold989 rf.registers\[26\]\[15\] VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ _2966_ _2980_ _2408_ _2990_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__o2bb2a_4
XANTENNA__5546__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8004_ _3126_ net580 _3963_ VGND VGND VPWR VPWR _3970_ sky130_fd_sc_hd__mux2_1
X_5216_ _1970_ _1971_ _1889_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6196_ _2895_ _2924_ _2363_ VGND VGND VPWR VPWR _2925_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5147_ _1766_ _1902_ _1672_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_86_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5078_ rf.registers\[4\]\[19\] rf.registers\[5\]\[19\] rf.registers\[6\]\[19\] rf.registers\[7\]\[19\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__mux4_1
XANTENNA__7379__A _3627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6283__A _3006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8906_ clknet_leaf_7_clk _0066_ VGND VGND VPWR VPWR rf.registers\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8837_ clknet_leaf_51_clk _1021_ VGND VGND VPWR VPWR rf.registers\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4809__S0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8768_ clknet_leaf_70_clk _0952_ VGND VGND VPWR VPWR rf.registers\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5482__S0 _1782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7719_ _3807_ VGND VGND VPWR VPWR _3819_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_117_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8699_ clknet_leaf_21_clk _0883_ VGND VGND VPWR VPWR rf.registers\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4531__A _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_152_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4677__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5537__S1 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5362__A _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7289__A _3590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4276__S1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7228__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4441__A _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5225__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold208 rf.registers\[31\]\[14\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold219 rf.registers\[10\]\[29\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4380_ rf.registers\[8\]\[1\] rf.registers\[9\]\[1\] rf.registers\[10\]\[1\] rf.registers\[11\]\[1\]
+ net117 _1053_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__mux4_1
XANTENNA__5064__A1_N _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6050_ _2785_ _2774_ _2786_ VGND VGND VPWR VPWR _2787_ sky130_fd_sc_hd__a21oi_1
X_5001_ _1669_ _1732_ _1756_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_147_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6952_ net223 _3130_ _3387_ VGND VGND VPWR VPWR _3396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5903_ _2567_ VGND VGND VPWR VPWR _2648_ sky130_fd_sc_hd__inv_2
X_6883_ _3359_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ _2581_ VGND VGND VPWR VPWR _2582_ sky130_fd_sc_hd__inv_2
X_8622_ clknet_leaf_41_clk _0806_ VGND VGND VPWR VPWR rf.registers\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5765_ _2323_ _2515_ VGND VGND VPWR VPWR _2516_ sky130_fd_sc_hd__and2_1
X_8553_ _4260_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7138__S _3498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7504_ _3705_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4351__A _1034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4716_ rf.registers\[8\]\[13\] rf.registers\[9\]\[13\] rf.registers\[10\]\[13\] rf.registers\[11\]\[13\]
+ _1291_ _1194_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4592__A1 _1171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8484_ _4224_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__clkbuf_1
X_5696_ net82 _1660_ VGND VGND VPWR VPWR _2450_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7435_ _3031_ net804 _3664_ VGND VGND VPWR VPWR _3669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6977__S _3375_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4647_ rf.registers\[28\]\[7\] rf.registers\[29\]\[7\] rf.registers\[30\]\[7\] rf.registers\[31\]\[7\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout2 _1172_ VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_96_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7366_ _3632_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
Xhold720 rf.registers\[8\]\[22\] VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold731 rf.registers\[6\]\[7\] VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
X_4578_ _1171_ _1323_ _1333_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__a21o_4
XFILLER_0_102_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold742 rf.registers\[10\]\[28\] VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold753 rf.registers\[16\]\[2\] VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__dlygate4sd3_1
X_6317_ net40 VGND VGND VPWR VPWR _3031_ sky130_fd_sc_hd__clkbuf_2
Xhold764 rf.registers\[21\]\[6\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd3_1
X_9105_ clknet_leaf_40_clk _0265_ VGND VGND VPWR VPWR rf.registers\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4497__S _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6278__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7297_ _3595_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
Xhold775 rf.registers\[14\]\[2\] VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5519__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold786 rf.registers\[25\]\[12\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 rf.registers\[27\]\[2\] VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd3_1
X_9036_ clknet_leaf_46_clk _0196_ VGND VGND VPWR VPWR rf.registers\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6248_ _2969_ _2973_ _2530_ VGND VGND VPWR VPWR _2974_ sky130_fd_sc_hd__mux2_1
X_6179_ _2017_ _1998_ VGND VGND VPWR VPWR _2909_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6217__S _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8432__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clone27_A _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7048__S _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5357__A _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5207__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6188__A _1978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7511__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold80 rf.registers\[7\]\[9\] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 rf.registers\[4\]\[9\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9251__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4436__A _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_63_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5446__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5550_ _1842_ _2305_ VGND VGND VPWR VPWR _2306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4501_ rf.registers\[20\]\[21\] rf.registers\[21\]\[21\] rf.registers\[22\]\[21\]
+ rf.registers\[23\]\[21\] _1220_ _1222_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__mux4_1
XANTENNA__6797__S _3304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5481_ _2233_ _2236_ _1828_ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4326__A1 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7220_ _3552_ _3553_ VGND VGND VPWR VPWR _3554_ sky130_fd_sc_hd__nand2_4
X_4432_ _1179_ _1186_ _1187_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__mux2_4
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4421__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7151_ _3516_ VGND VGND VPWR VPWR _3517_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4363_ rf.registers\[0\]\[2\] rf.registers\[1\]\[2\] rf.registers\[2\]\[2\] rf.registers\[3\]\[2\]
+ net94 _1061_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6102_ _1512_ _2835_ net1160 _2658_ _2536_ VGND VGND VPWR VPWR _2836_ sky130_fd_sc_hd__a41o_1
XFILLER_0_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7082_ net44 VGND VGND VPWR VPWR _3472_ sky130_fd_sc_hd__buf_2
X_4294_ net7 VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__clkinv_4
XANTENNA__5826__A1 _2105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _2770_ VGND VGND VPWR VPWR _2771_ sky130_fd_sc_hd__inv_2
XANTENNA__7421__S _3627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5730__A _2080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer23 net104 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
XANTENNA__4346__A _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer34 _1542_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7984_ _3959_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer45 _1166_ VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_107_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4488__S1 _1208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6935_ _3375_ VGND VGND VPWR VPWR _3387_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8252__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
X_6866_ _3350_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8605_ clknet_leaf_15_clk _0789_ VGND VGND VPWR VPWR rf.registers\[22\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6280__B net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5817_ _2565_ VGND VGND VPWR VPWR _2566_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6797_ net234 _3111_ _3304_ VGND VGND VPWR VPWR _3314_ sky130_fd_sc_hd__mux2_1
X_9585_ clknet_leaf_29_clk _0745_ VGND VGND VPWR VPWR rf.registers\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8536_ _4251_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__clkbuf_1
X_5748_ _2418_ _2499_ _1147_ VGND VGND VPWR VPWR _2500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8467_ _4215_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__clkbuf_1
X_5679_ _2307_ _2325_ _1148_ VGND VGND VPWR VPWR _2433_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_3_5__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5514__B1 _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7418_ _3659_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__clkbuf_1
X_8398_ net785 _3474_ _4169_ VGND VGND VPWR VPWR _4179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold550 rf.registers\[29\]\[1\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__dlygate4sd3_1
X_7349_ _3622_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
Xhold561 rf.registers\[8\]\[17\] VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 rf.registers\[19\]\[15\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5116__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold583 rf.registers\[29\]\[27\] VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 rf.registers\[27\]\[1\] VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9274__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9019_ clknet_leaf_34_clk _0179_ VGND VGND VPWR VPWR rf.registers\[31\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5640__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5045__A2 _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8162__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5428__S0 _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5753__B1 _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4651__S1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4403__S1 _1028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput70 net70 VGND VGND VPWR VPWR alu_out[29] sky130_fd_sc_hd__buf_6
XFILLER_0_37_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output65_A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4865__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8337__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5550__A _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6233__A1 _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4981_ rf.registers\[16\]\[22\] rf.registers\[17\]\[22\] rf.registers\[18\]\[22\]
+ rf.registers\[19\]\[22\] _1734_ _1735_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6720_ _3033_ net1028 _3267_ VGND VGND VPWR VPWR _3273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6651_ _3236_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5602_ net82 _2287_ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6582_ _3031_ net1086 _3195_ VGND VGND VPWR VPWR _3200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9370_ clknet_leaf_37_clk _0530_ VGND VGND VPWR VPWR rf.registers\[20\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8321_ _4138_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__clkbuf_1
X_5533_ _1169_ _2272_ _2288_ VGND VGND VPWR VPWR _2289_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8252_ _3101_ net1004 _4097_ VGND VGND VPWR VPWR _4102_ sky130_fd_sc_hd__mux2_1
X_5464_ _2216_ _2219_ _1699_ VGND VGND VPWR VPWR _2220_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7203_ _3544_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
X_4415_ _1170_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__buf_8
XFILLER_0_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8183_ _4065_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__clkbuf_1
X_5395_ _2147_ _2150_ net4 VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7134_ _3507_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
X_4346_ _1071_ _1101_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7065_ net411 _3460_ _3456_ VGND VGND VPWR VPWR _3461_ sky130_fd_sc_hd__mux2_1
X_4277_ rf.registers\[24\]\[4\] rf.registers\[25\]\[4\] rf.registers\[26\]\[4\] rf.registers\[27\]\[4\]
+ _1027_ _1029_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__mux4_1
X_6016_ _2496_ _2754_ VGND VGND VPWR VPWR _2755_ sky130_fd_sc_hd__and2_1
XANTENNA__5680__C1 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6990__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7967_ net254 _3452_ _3915_ VGND VGND VPWR VPWR _3950_ sky130_fd_sc_hd__mux2_1
XANTENNA__5432__C1 _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _3378_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_120_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7898_ _3913_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6849_ net211 _3095_ _3340_ VGND VGND VPWR VPWR _3342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9568_ clknet_leaf_70_clk _0728_ VGND VGND VPWR VPWR rf.registers\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4633__S1 _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8519_ _4242_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__clkbuf_1
X_9499_ clknet_leaf_34_clk _0659_ VGND VGND VPWR VPWR rf.registers\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold380 rf.registers\[3\]\[17\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 rf.registers\[17\]\[5\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7996__S _3963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7963__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_25_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4624__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer3 net84 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7236__S _3555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7479__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_39_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5180_ rf.registers\[0\]\[29\] rf.registers\[1\]\[29\] rf.registers\[2\]\[29\] rf.registers\[3\]\[29\]
+ _1895_ _1897_ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__mux4_1
XANTENNA__8067__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6376__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8870_ clknet_leaf_72_clk _0030_ VGND VGND VPWR VPWR rf.registers\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7821_ net358 _3442_ _3866_ VGND VGND VPWR VPWR _3873_ sky130_fd_sc_hd__mux2_1
XANTENNA__6315__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4312__S0 _1065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4964_ _1719_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__buf_4
X_7752_ _3836_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_16_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
X_6703_ _3263_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4895_ rf.registers\[8\]\[0\] rf.registers\[9\]\[0\] rf.registers\[10\]\[0\] rf.registers\[11\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7683_ net615 _3508_ _3794_ VGND VGND VPWR VPWR _3800_ sky130_fd_sc_hd__mux2_1
X_9422_ clknet_leaf_29_clk _0582_ VGND VGND VPWR VPWR rf.registers\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6634_ _3083_ net814 _3217_ VGND VGND VPWR VPWR _3227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9353_ clknet_leaf_51_clk _0513_ VGND VGND VPWR VPWR rf.registers\[20\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6565_ _3189_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7146__S _3455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5455__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8304_ _3013_ net1144 _4119_ VGND VGND VPWR VPWR _4129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5516_ _1638_ _2271_ VGND VGND VPWR VPWR _2272_ sky130_fd_sc_hd__or2_1
X_9284_ clknet_leaf_47_clk _0444_ VGND VGND VPWR VPWR rf.registers\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6496_ _3151_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8131__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5447_ rf.registers\[12\]\[10\] rf.registers\[13\]\[10\] rf.registers\[14\]\[10\]
+ rf.registers\[15\]\[10\] _2117_ _2118_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__mux4_1
X_8235_ _4092_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5378_ _2132_ _2133_ _1711_ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__mux2_1
X_8166_ net844 _3446_ _4047_ VGND VGND VPWR VPWR _4056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4329_ net47 _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__nor2_2
X_7117_ net388 _3495_ _3477_ VGND VGND VPWR VPWR _3496_ sky130_fd_sc_hd__mux2_1
X_8097_ _4019_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__clkbuf_1
X_7048_ net490 _3448_ _3435_ VGND VGND VPWR VPWR _3449_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4551__S0 net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8999_ clknet_leaf_66_clk _0159_ VGND VGND VPWR VPWR rf.registers\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7945__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4534__A _1065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5420__A2 _2175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4854__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8440__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8370__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8122__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6895__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5031__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6684__A1 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4790__S0 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5304__S _1685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4998__A1 _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7936__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__S1 _1823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4444__A _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4680_ _1434_ _1435_ _1178_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6350_ _3053_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5301_ _1828_ _2056_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6281_ net9 _3004_ VGND VGND VPWR VPWR _3005_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_73_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5232_ rf.registers\[12\]\[26\] rf.registers\[13\]\[26\] rf.registers\[14\]\[26\]
+ rf.registers\[15\]\[26\] _1896_ _1898_ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__mux4_1
XANTENNA__6675__A1 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8020_ _3978_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_5_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__5883__C1 _2504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5163_ _1823_ VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__clkbuf_4
X_5094_ rf.registers\[8\]\[17\] rf.registers\[9\]\[17\] rf.registers\[10\]\[17\] rf.registers\[11\]\[17\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8922_ clknet_leaf_17_clk _0082_ VGND VGND VPWR VPWR rf.registers\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8525__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8853_ clknet_leaf_32_clk _0013_ VGND VGND VPWR VPWR rf.registers\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7804_ net170 _3493_ _3855_ VGND VGND VPWR VPWR _3864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8784_ clknet_leaf_12_clk _0968_ VGND VGND VPWR VPWR rf.registers\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_5996_ _2733_ _2735_ _1879_ VGND VGND VPWR VPWR _2736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4836__S1 _1078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7735_ _3827_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__clkbuf_1
X_4947_ _1702_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__8260__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7666_ net540 _3491_ _3783_ VGND VGND VPWR VPWR _3791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4878_ _1239_ _1625_ _1629_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__a2bb2o_2
X_9405_ clknet_leaf_15_clk _0565_ VGND VGND VPWR VPWR rf.registers\[24\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5166__A1 _1766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6617_ _3218_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7597_ _3754_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_65_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9336_ clknet_leaf_26_clk _0496_ VGND VGND VPWR VPWR rf.registers\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6548_ net422 _3137_ _3179_ VGND VGND VPWR VPWR _3181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9267_ clknet_leaf_35_clk _0427_ VGND VGND VPWR VPWR rf.registers\[23\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6479_ net1054 _3141_ _3135_ VGND VGND VPWR VPWR _3142_ sky130_fd_sc_hd__mux2_1
XANTENNA__5013__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8218_ net419 _3497_ _4083_ VGND VGND VPWR VPWR _4084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9198_ clknet_leaf_44_clk _0358_ VGND VGND VPWR VPWR rf.registers\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8149_ _4024_ VGND VGND VPWR VPWR _4047_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__6107__B_N _1779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7615__A0 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4524__S0 net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4827__S1 _1183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8170__S _4024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8343__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5252__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5004__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4439__A _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8345__S _4144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8031__A0 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5850_ _2229_ _2597_ VGND VGND VPWR VPWR _2598_ sky130_fd_sc_hd__xor2_2
XFILLER_0_76_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4801_ _1088_ _1556_ net8 VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_66_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4818__S1 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5781_ _2255_ _2355_ _2364_ _2337_ VGND VGND VPWR VPWR _2532_ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7520_ _3048_ net699 _3711_ VGND VGND VPWR VPWR _3714_ sky130_fd_sc_hd__mux2_1
X_4732_ rf.registers\[0\]\[14\] rf.registers\[1\]\[14\] rf.registers\[2\]\[14\] rf.registers\[3\]\[14\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7451_ _3677_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__clkbuf_1
X_4663_ rf.registers\[16\]\[23\] rf.registers\[17\]\[23\] rf.registers\[18\]\[23\]
+ rf.registers\[19\]\[23\] _1351_ _1352_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5209__S _1745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6402_ _3088_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7382_ _3046_ net1142 _3639_ VGND VGND VPWR VPWR _3641_ sky130_fd_sc_hd__mux2_1
X_4594_ _1238_ _1278_ _1316_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__or4_4
Xhold902 rf.registers\[1\]\[27\] VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold913 rf.registers\[13\]\[21\] VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__dlygate4sd3_1
X_9121_ clknet_leaf_57_clk _0281_ VGND VGND VPWR VPWR rf.registers\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6333_ _3041_ net843 _3023_ VGND VGND VPWR VPWR _3042_ sky130_fd_sc_hd__mux2_1
Xhold924 rf.registers\[28\]\[20\] VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 rf.registers\[24\]\[1\] VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold946 rf.registers\[14\]\[5\] VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6648__A1 _3099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7845__A0 _3103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold957 rf.registers\[30\]\[18\] VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 rf.registers\[23\]\[12\] VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__dlygate4sd3_1
X_6264_ _2988_ _2989_ VGND VGND VPWR VPWR _2990_ sky130_fd_sc_hd__nor2_1
X_9052_ clknet_leaf_16_clk _0212_ VGND VGND VPWR VPWR rf.registers\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold979 rf.registers\[29\]\[31\] VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__dlygate4sd3_1
X_8003_ _3969_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__clkbuf_1
X_5215_ rf.registers\[12\]\[27\] rf.registers\[13\]\[27\] rf.registers\[14\]\[27\]
+ rf.registers\[15\]\[27\] _1918_ _1919_ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__mux4_1
XANTENNA__4349__A _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6195_ _2923_ _2384_ VGND VGND VPWR VPWR _2924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5146_ _1899_ _1900_ _1901_ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5077_ _1700_ _1832_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__nand2_1
XANTENNA__5084__B1 _1839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8905_ clknet_leaf_45_clk _0065_ VGND VGND VPWR VPWR rf.registers\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8836_ clknet_leaf_51_clk _1020_ VGND VGND VPWR VPWR rf.registers\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4809__S1 _1053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5387__A1 _1169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8767_ clknet_leaf_71_clk _0951_ VGND VGND VPWR VPWR rf.registers\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_5979_ _2569_ _2719_ _2104_ VGND VGND VPWR VPWR _2720_ sky130_fd_sc_hd__mux2_1
XANTENNA__5908__A _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5482__S1 _1680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7718_ _3818_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8698_ clknet_leaf_18_clk _0882_ VGND VGND VPWR VPWR rf.registers\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7649_ net753 _3474_ _3772_ VGND VGND VPWR VPWR _3782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9319_ clknet_leaf_65_clk _0479_ VGND VGND VPWR VPWR rf.registers\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4958__S _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7334__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8013__A0 _3134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8564__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7509__S _3700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5029__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5225__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold209 rf.registers\[17\]\[16\] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4868__S _1259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4353__A2 _1088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5000_ _1668_ _1755_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8252__A0 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8075__S _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6802__A1 _3116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6951_ _3395_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5161__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8004__A0 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5902_ _2644_ _2646_ VGND VGND VPWR VPWR _2647_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6882_ net384 _3128_ _3351_ VGND VGND VPWR VPWR _3359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8621_ clknet_leaf_41_clk _0805_ VGND VGND VPWR VPWR rf.registers\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5833_ _2230_ _2580_ _1839_ VGND VGND VPWR VPWR _2581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5728__A _2062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7419__S _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8552_ net705 net23 _4255_ VGND VGND VPWR VPWR _4260_ sky130_fd_sc_hd__mux2_1
XANTENNA__4577__C1 _1215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5764_ _1083_ _2514_ VGND VGND VPWR VPWR _2515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7503_ _3031_ net1134 _3700_ VGND VGND VPWR VPWR _3705_ sky130_fd_sc_hd__mux2_1
X_4715_ _1467_ _1470_ _1071_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8483_ net725 net22 _4216_ VGND VGND VPWR VPWR _4224_ sky130_fd_sc_hd__mux2_1
X_5695_ _2080_ _2448_ VGND VGND VPWR VPWR _2449_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7434_ _3668_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4646_ _1400_ _1401_ _1107_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold710 rf.registers\[11\]\[15\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7365_ _3029_ net1108 _3628_ VGND VGND VPWR VPWR _3632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4577_ _1327_ _1329_ _1332_ _1187_ _1215_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__o221a_1
Xhold721 rf.registers\[0\]\[31\] VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7154__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold732 rf.registers\[15\]\[29\] VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold743 rf.registers\[24\]\[2\] VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd3_1
X_9104_ clknet_leaf_3_clk _0264_ VGND VGND VPWR VPWR rf.registers\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6316_ _3030_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold754 rf.registers\[26\]\[1\] VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold765 rf.registers\[11\]\[18\] VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlygate4sd3_1
X_7296_ _3029_ net806 _3591_ VGND VGND VPWR VPWR _3595_ sky130_fd_sc_hd__mux2_1
Xhold776 rf.registers\[19\]\[28\] VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 rf.registers\[25\]\[18\] VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd3_1
X_9035_ clknet_leaf_2_clk _0195_ VGND VGND VPWR VPWR rf.registers\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold798 rf.registers\[26\]\[17\] VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4727__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6247_ _2972_ VGND VGND VPWR VPWR _2973_ sky130_fd_sc_hd__inv_2
X_6178_ _2444_ _2864_ VGND VGND VPWR VPWR _2908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5129_ rf.registers\[24\]\[31\] rf.registers\[25\]\[31\] rf.registers\[26\]\[31\]
+ rf.registers\[27\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_127_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5402__S net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6254__C1 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8546__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8819_ clknet_leaf_33_clk _1003_ VGND VGND VPWR VPWR rf.registers\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7329__S _3602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5207__S1 _1768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4688__S _1211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6469__A _3092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6408__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold70 rf.registers\[17\]\[12\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 rf.registers\[9\]\[25\] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 rf.registers\[14\]\[11\] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5143__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8537__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5446__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4452__A _1174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4500_ _1246_ _1239_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__o21ai_4
X_5480_ _2234_ _2235_ _1685_ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4431_ _1071_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6379__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4362_ _1107_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__or2_1
X_7150_ _3411_ _3302_ VGND VGND VPWR VPWR _3516_ sky130_fd_sc_hd__nor2_4
XFILLER_0_67_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6101_ net104 net133 VGND VGND VPWR VPWR _2835_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7081_ _3471_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
X_4293_ rf.registers\[0\]\[4\] rf.registers\[1\]\[4\] rf.registers\[2\]\[4\] rf.registers\[3\]\[4\]
+ net103 _1044_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__mux4_1
XANTENNA__4709__S0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6032_ _2744_ _2763_ VGND VGND VPWR VPWR _2770_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7028__A1 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6318__S _3023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer13 _2506_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer24 _1298_ VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__5134__S0 _1889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7983_ _3105_ net846 _3952_ VGND VGND VPWR VPWR _3959_ sky130_fd_sc_hd__mux2_1
Xrebuffer35 _2711_ VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer46 _1166_ VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_89_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8533__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6934_ _3386_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6865_ net145 _3111_ _3340_ VGND VGND VPWR VPWR _3350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7200__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8604_ clknet_leaf_16_clk _0788_ VGND VGND VPWR VPWR rf.registers\[22\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4362__A _1107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5816_ _2361_ _2357_ VGND VGND VPWR VPWR _2565_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9584_ clknet_leaf_12_clk _0744_ VGND VGND VPWR VPWR rf.registers\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6796_ _3313_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_98_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6988__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8535_ net347 net15 _4244_ VGND VGND VPWR VPWR _4251_ sky130_fd_sc_hd__mux2_1
X_5747_ _2498_ VGND VGND VPWR VPWR _2499_ sky130_fd_sc_hd__inv_2
XANTENNA__5762__B2 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8466_ net521 net45 _4205_ VGND VGND VPWR VPWR _4215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5678_ _2083_ VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__inv_2
XANTENNA__5514__A1 _1828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7417_ _3081_ net837 _3650_ VGND VGND VPWR VPWR _3659_ sky130_fd_sc_hd__mux2_1
X_4629_ _1370_ _1384_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__nand2_1
X_8397_ _4178_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold540 rf.registers\[16\]\[17\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold551 rf.registers\[15\]\[18\] VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
X_7348_ _3081_ net742 _3613_ VGND VGND VPWR VPWR _3622_ sky130_fd_sc_hd__mux2_1
Xhold562 rf.registers\[0\]\[12\] VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 rf.registers\[23\]\[15\] VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold584 rf.registers\[27\]\[8\] VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold595 rf.registers\[28\]\[28\] VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7279_ _3585_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_9018_ clknet_leaf_35_clk _0178_ VGND VGND VPWR VPWR rf.registers\[31\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5373__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4971__S _1726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7059__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5368__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5428__S1 _1716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5202__B1 _1957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7583__A _3735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput60 net60 VGND VGND VPWR VPWR alu_out[1] sky130_fd_sc_hd__buf_6
Xoutput71 net71 VGND VGND VPWR VPWR alu_out[2] sky130_fd_sc_hd__buf_4
XANTENNA__7522__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5364__S0 _2117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5550__B _2305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output58_A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6662__A _3230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4980_ rf.registers\[20\]\[22\] rf.registers\[21\]\[22\] rf.registers\[22\]\[22\]
+ rf.registers\[23\]\[22\] _1734_ _1735_ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5278__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6650_ net629 _3101_ _3231_ VGND VGND VPWR VPWR _3236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5601_ _2348_ _2355_ _1879_ VGND VGND VPWR VPWR _2356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6581_ _3199_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8320_ net157 _3464_ _4133_ VGND VGND VPWR VPWR _4138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6601__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5532_ _1800_ _2287_ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__nor2_1
X_8251_ _4101_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5463_ _2217_ _2218_ _1685_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7202_ net827 _3506_ _3539_ VGND VGND VPWR VPWR _3544_ sky130_fd_sc_hd__mux2_1
X_4414_ _1057_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__buf_4
X_8182_ net523 _3462_ _4061_ VGND VGND VPWR VPWR _4065_ sky130_fd_sc_hd__mux2_1
X_5394_ _2148_ _2149_ _1684_ VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7133_ net543 _3506_ _3498_ VGND VGND VPWR VPWR _3507_ sky130_fd_sc_hd__mux2_1
X_4345_ _1099_ _1100_ _1048_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7064_ net36 VGND VGND VPWR VPWR _3460_ sky130_fd_sc_hd__buf_2
X_4276_ rf.registers\[28\]\[4\] rf.registers\[29\]\[4\] rf.registers\[30\]\[4\] rf.registers\[31\]\[4\]
+ _1027_ _1029_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__mux4_1
XANTENNA__5355__S0 _1703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6015_ _2751_ _2753_ _2252_ VGND VGND VPWR VPWR _2754_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5107__S0 _1705_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _3949_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6917_ net597 _3095_ _3376_ VGND VGND VPWR VPWR _3378_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4786__A2 _1025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7897_ _3015_ net673 _3879_ VGND VGND VPWR VPWR _3913_ sky130_fd_sc_hd__mux2_1
XANTENNA__5188__A _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6848_ _3341_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9567_ clknet_leaf_71_clk _0727_ VGND VGND VPWR VPWR rf.registers\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6779_ net272 _3089_ _3304_ VGND VGND VPWR VPWR _3305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7607__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8518_ net349 net36 _3007_ VGND VGND VPWR VPWR _4242_ sky130_fd_sc_hd__mux2_1
X_9498_ clknet_leaf_37_clk _0658_ VGND VGND VPWR VPWR rf.registers\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8449_ _4206_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold370 rf.registers\[24\]\[7\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8438__S _4191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold381 rf.registers\[26\]\[0\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7342__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold392 rf.registers\[26\]\[13\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7660__A1 _3485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1070 rf.registers\[30\]\[19\] VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5974__B2 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer4 net85 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_58_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4876__S _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5337__S0 _1641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5662__B1 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7820_ _3872_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4905__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7751_ _3075_ net808 _3830_ VGND VGND VPWR VPWR _3836_ sky130_fd_sc_hd__mux2_1
XANTENNA__4312__S1 _1066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4963_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6702_ net245 _3013_ _3253_ VGND VGND VPWR VPWR _3263_ sky130_fd_sc_hd__mux2_1
X_7682_ _3799_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__clkbuf_1
X_4894_ _1646_ _1649_ net4 VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__mux2_1
XANTENNA__5980__A4 _2472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9421_ clknet_leaf_44_clk _0581_ VGND VGND VPWR VPWR rf.registers\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6633_ _3226_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7427__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9352_ clknet_leaf_48_clk _0512_ VGND VGND VPWR VPWR rf.registers\[20\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6564_ net737 _3013_ _3179_ VGND VGND VPWR VPWR _3189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8303_ _4128_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5515_ _1670_ _2262_ _2266_ _2270_ VGND VGND VPWR VPWR _2271_ sky130_fd_sc_hd__a2bb2o_1
X_9283_ clknet_leaf_68_clk _0443_ VGND VGND VPWR VPWR rf.registers\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6495_ net906 _3015_ _3092_ VGND VGND VPWR VPWR _3151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8234_ net195 _3446_ _4083_ VGND VGND VPWR VPWR _4092_ sky130_fd_sc_hd__mux2_1
X_5446_ rf.registers\[8\]\[10\] rf.registers\[9\]\[10\] rf.registers\[10\]\[10\] rf.registers\[11\]\[10\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8258__S _4097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8165_ _4055_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__clkbuf_1
X_5377_ rf.registers\[12\]\[14\] rf.registers\[13\]\[14\] rf.registers\[14\]\[14\]
+ rf.registers\[15\]\[14\] _2113_ _2114_ VGND VGND VPWR VPWR _2133_ sky130_fd_sc_hd__mux4_1
XANTENNA__7162__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7116_ net24 VGND VGND VPWR VPWR _3495_ sky130_fd_sc_hd__buf_2
XANTENNA__5328__S0 _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4328_ net48 _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__nand2_1
X_8096_ net317 _3444_ _4011_ VGND VGND VPWR VPWR _4019_ sky130_fd_sc_hd__mux2_1
X_7047_ net35 VGND VGND VPWR VPWR _3448_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4551__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6506__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8998_ clknet_leaf_0_clk _0158_ VGND VGND VPWR VPWR rf.registers\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5405__B1 _1800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5500__S0 _1733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7949_ net978 _3502_ _3938_ VGND VGND VPWR VPWR _3941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5646__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8168__S _4047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4790__S1 _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5644__B1 _1799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7800__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7101__A net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7247__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5300_ _2054_ _2055_ _1712_ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7321__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6280_ net10 net46 VGND VGND VPWR VPWR _3004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5231_ _1983_ _1986_ _1766_ VGND VGND VPWR VPWR _1987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5162_ _1822_ VGND VGND VPWR VPWR _1918_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5093_ _1845_ _1848_ _1697_ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__mux2_1
X_8921_ clknet_leaf_20_clk _0081_ VGND VGND VPWR VPWR rf.registers\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_3_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7388__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8852_ clknet_leaf_30_clk _0012_ VGND VGND VPWR VPWR rf.registers\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8107__A _4024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5230__S _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7803_ _3863_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5938__A1 _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8783_ clknet_leaf_28_clk _0967_ VGND VGND VPWR VPWR rf.registers\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5995_ _2703_ _2734_ _2347_ VGND VGND VPWR VPWR _2735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8541__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7734_ _3058_ net823 _3819_ VGND VGND VPWR VPWR _3827_ sky130_fd_sc_hd__mux2_1
X_4946_ _1701_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7665_ _3790_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _1254_ _1632_ _1170_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9404_ clknet_leaf_17_clk _0564_ VGND VGND VPWR VPWR rf.registers\[24\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6616_ _3064_ net486 _3217_ VGND VGND VPWR VPWR _3218_ sky130_fd_sc_hd__mux2_1
X_7596_ _3056_ net907 _3747_ VGND VGND VPWR VPWR _3754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9335_ clknet_leaf_33_clk _0495_ VGND VGND VPWR VPWR rf.registers\[21\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6996__S _3413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6547_ _3180_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9266_ clknet_leaf_38_clk _0426_ VGND VGND VPWR VPWR rf.registers\[23\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6478_ net29 VGND VGND VPWR VPWR _3141_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8217_ _4060_ VGND VGND VPWR VPWR _4083_ sky130_fd_sc_hd__buf_4
XANTENNA__5323__C1 _1640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5429_ rf.registers\[12\]\[11\] rf.registers\[13\]\[11\] rf.registers\[14\]\[11\]
+ rf.registers\[15\]\[11\] _1704_ _1707_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9197_ clknet_leaf_49_clk _0357_ VGND VGND VPWR VPWR rf.registers\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8148_ _4046_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__clkbuf_1
X_8079_ net863 _3495_ _4000_ VGND VGND VPWR VPWR _4010_ sky130_fd_sc_hd__mux2_1
XANTENNA__4524__S1 _1279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4280__A _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5315__S net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6935__A _3375_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7530__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4455__A _1198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7766__A _3843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6042__B1 _2333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4800_ _1554_ _1555_ _1107_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _2403_ _2348_ _1879_ VGND VGND VPWR VPWR _2531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4731_ _1198_ _1486_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7450_ _3046_ net1090 _3675_ VGND VGND VPWR VPWR _3677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4662_ rf.registers\[28\]\[23\] rf.registers\[29\]\[23\] rf.registers\[30\]\[23\]
+ rf.registers\[31\]\[23\] _1267_ _1268_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6401_ _3087_ net601 _3022_ VGND VGND VPWR VPWR _3088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7381_ _3640_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4593_ _1334_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7705__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9120_ clknet_leaf_60_clk _0280_ VGND VGND VPWR VPWR rf.registers\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold903 rf.registers\[21\]\[2\] VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6332_ net45 VGND VGND VPWR VPWR _3041_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__8098__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold914 rf.registers\[15\]\[27\] VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 rf.registers\[31\]\[5\] VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold936 rf.registers\[26\]\[12\] VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 rf.registers\[28\]\[23\] VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 rf.registers\[30\]\[0\] VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__dlygate4sd3_1
X_9051_ clknet_leaf_36_clk _0211_ VGND VGND VPWR VPWR rf.registers\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold969 rf.registers\[29\]\[9\] VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__dlygate4sd3_1
X_6263_ _2952_ _2987_ _2986_ VGND VGND VPWR VPWR _2989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8002_ _3124_ net390 _3963_ VGND VGND VPWR VPWR _3969_ sky130_fd_sc_hd__mux2_1
X_5214_ rf.registers\[8\]\[27\] rf.registers\[9\]\[27\] rf.registers\[10\]\[27\] rf.registers\[11\]\[27\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__mux4_1
X_6194_ _1669_ _1997_ VGND VGND VPWR VPWR _2923_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5145_ _1726_ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5076_ _1830_ _1831_ _1686_ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__mux2_1
X_8904_ clknet_leaf_63_clk _0064_ VGND VGND VPWR VPWR rf.registers\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8835_ clknet_leaf_53_clk _1019_ VGND VGND VPWR VPWR rf.registers\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8271__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8766_ clknet_leaf_0_clk _0950_ VGND VGND VPWR VPWR rf.registers\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5978_ _2650_ _2718_ _2251_ VGND VGND VPWR VPWR _2719_ sky130_fd_sc_hd__mux2_1
X_7717_ _3041_ net693 _3808_ VGND VGND VPWR VPWR _3818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4929_ _1684_ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8697_ clknet_leaf_19_clk _0881_ VGND VGND VPWR VPWR rf.registers\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_7648_ _3781_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7579_ _3039_ net710 _3736_ VGND VGND VPWR VPWR _3745_ sky130_fd_sc_hd__mux2_1
XANTENNA__7615__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9318_ clknet_leaf_0_clk _0478_ VGND VGND VPWR VPWR rf.registers\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9249_ clknet_leaf_58_clk _0409_ VGND VGND VPWR VPWR rf.registers\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7350__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7524__A0 _3052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7827__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_84_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8356__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6950_ net855 _3128_ _3387_ VGND VGND VPWR VPWR _3395_ sky130_fd_sc_hd__mux2_1
XANTENNA__5161__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5901_ net112 _2636_ _2645_ VGND VGND VPWR VPWR _2646_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6881_ _3358_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8620_ clknet_leaf_50_clk _0804_ VGND VGND VPWR VPWR rf.registers\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_93_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5832_ _2287_ VGND VGND VPWR VPWR _2580_ sky130_fd_sc_hd__inv_2
XANTENNA__4913__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8551_ _4259_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__clkbuf_1
X_5763_ _1060_ net95 _2411_ VGND VGND VPWR VPWR _2514_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7502_ _3704_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
X_4714_ _1468_ _1469_ _1036_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8482_ _4223_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__clkbuf_1
X_5694_ net84 _2447_ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7433_ _3029_ net283 _3664_ VGND VGND VPWR VPWR _3668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4645_ rf.registers\[16\]\[7\] rf.registers\[17\]\[7\] rf.registers\[18\]\[7\] rf.registers\[19\]\[7\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__mux4_1
XANTENNA__4424__S0 _1173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7435__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold700 rf.registers\[13\]\[7\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7364_ _3631_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4576_ _1330_ _1331_ _1259_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold711 rf.registers\[22\]\[21\] VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold722 rf.registers\[25\]\[4\] VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold733 rf.registers\[3\]\[7\] VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
X_9103_ clknet_leaf_9_clk _0263_ VGND VGND VPWR VPWR rf.registers\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6315_ _3029_ net840 _3023_ VGND VGND VPWR VPWR _3030_ sky130_fd_sc_hd__mux2_1
Xhold744 rf.registers\[21\]\[31\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 rf.registers\[26\]\[28\] VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__dlygate4sd3_1
X_7295_ _3594_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
Xhold766 rf.registers\[13\]\[2\] VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 rf.registers\[23\]\[5\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd3_1
X_9034_ clknet_leaf_8_clk _0194_ VGND VGND VPWR VPWR rf.registers\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold788 rf.registers\[1\]\[22\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 rf.registers\[30\]\[8\] VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _2970_ _2971_ _1126_ VGND VGND VPWR VPWR _2972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4727__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6177_ _2626_ _2797_ VGND VGND VPWR VPWR _2907_ sky130_fd_sc_hd__nor2_1
XANTENNA__7170__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5128_ _1883_ VGND VGND VPWR VPWR _1884_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ _1700_ _1814_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_48_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6514__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8818_ clknet_leaf_25_clk _1002_ VGND VGND VPWR VPWR rf.registers\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8749_ clknet_leaf_8_clk _0933_ VGND VGND VPWR VPWR rf.registers\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4663__S0 _1351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7809__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8176__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7080__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8234__A1 _3446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold60 rf.registers\[5\]\[11\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 rf.registers\[9\]\[23\] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 rf.registers\[18\]\[13\] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 rf.registers\[12\]\[14\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5143__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6548__A1 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4406__S0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7255__S _3566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4430_ _1180_ _1185_ _1178_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__mux2_1
XANTENNA_2 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4361_ rf.registers\[4\]\[2\] rf.registers\[5\]\[2\] rf.registers\[6\]\[2\] rf.registers\[7\]\[2\]
+ net101 _1066_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6100_ _2496_ _2822_ _2826_ _2834_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__a211o_1
X_7080_ net815 _3470_ _3456_ VGND VGND VPWR VPWR _3471_ sky130_fd_sc_hd__mux2_1
XANTENNA__8473__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4292_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__buf_4
XANTENNA__4709__S1 _1029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6031_ _1820_ _2768_ VGND VGND VPWR VPWR _2769_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_91_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8086__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4908__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer14 _1573_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd1_1
X_7982_ _3958_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6787__A1 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5134__S1 _1773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer36 _1399_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer47 _2664_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd1_1
X_6933_ net173 _3111_ _3376_ VGND VGND VPWR VPWR _3386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6864_ _3349_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7736__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5815_ _2561_ _2563_ VGND VGND VPWR VPWR _2564_ sky130_fd_sc_hd__xnor2_1
X_8603_ clknet_leaf_34_clk _0787_ VGND VGND VPWR VPWR rf.registers\[22\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_9583_ clknet_leaf_27_clk _0743_ VGND VGND VPWR VPWR rf.registers\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6795_ net197 _3109_ _3304_ VGND VGND VPWR VPWR _3313_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4645__S0 _1104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8534_ _4250_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5746_ _2064_ _2307_ VGND VGND VPWR VPWR _2498_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_98_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4789__S _1034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8465_ _4214_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__clkbuf_1
X_5677_ _2430_ _2289_ _2363_ VGND VGND VPWR VPWR _2431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5474__A _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7416_ _3658_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4628_ _1171_ _1375_ _1379_ _1383_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8396_ net252 _3472_ _4169_ VGND VGND VPWR VPWR _4178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5070__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold530 rf.registers\[8\]\[25\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7347_ _3621_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
Xhold541 rf.registers\[11\]\[1\] VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _1171_ _1306_ _1310_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__o2bb2a_4
Xhold552 rf.registers\[0\]\[5\] VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 rf.registers\[17\]\[29\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 rf.registers\[9\]\[16\] VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8464__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold585 rf.registers\[19\]\[11\] VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__dlygate4sd3_1
X_7278_ _3079_ net665 _3577_ VGND VGND VPWR VPWR _3585_ sky130_fd_sc_hd__mux2_1
Xhold596 rf.registers\[29\]\[28\] VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9017_ clknet_leaf_19_clk _0177_ VGND VGND VPWR VPWR rf.registers\[31\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6229_ _2953_ _2954_ VGND VGND VPWR VPWR _2956_ sky130_fd_sc_hd__nand2_1
XANTENNA__5413__S _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5373__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5202__A1 _1777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4699__S _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6702__A1 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5061__S0 _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput50 net50 VGND VGND VPWR VPWR alu_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_102_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput61 net61 VGND VGND VPWR VPWR alu_out[20] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VGND VGND VPWR VPWR alu_out[30] sky130_fd_sc_hd__buf_8
XANTENNA__5364__S1 _2118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7104__A net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8207__A1 _3487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4875__S0 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4463__A _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5278__B _2033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7194__A1 _3497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5600_ _2351_ _2354_ _2347_ VGND VGND VPWR VPWR _2355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6580_ _3029_ net999 _3195_ VGND VGND VPWR VPWR _3199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5531_ net1163 _2286_ VGND VGND VPWR VPWR _2287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5294__A _1673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8250_ _3099_ net387 _4097_ VGND VGND VPWR VPWR _4101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5462_ rf.registers\[24\]\[8\] rf.registers\[25\]\[8\] rf.registers\[26\]\[8\] rf.registers\[27\]\[8\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5052__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7201_ _3543_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
X_4413_ _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8181_ _4064_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5393_ rf.registers\[24\]\[13\] rf.registers\[25\]\[13\] rf.registers\[26\]\[13\]
+ rf.registers\[27\]\[13\] _1673_ _1690_ VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__mux4_1
XANTENNA__7713__S _3808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7132_ net30 VGND VGND VPWR VPWR _3506_ sky130_fd_sc_hd__buf_2
X_4344_ rf.registers\[12\]\[3\] rf.registers\[13\]\[3\] rf.registers\[14\]\[3\] rf.registers\[15\]\[3\]
+ net103 _1044_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7063_ _3459_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
X_4275_ rf.registers\[16\]\[4\] rf.registers\[17\]\[4\] rf.registers\[18\]\[4\] rf.registers\[19\]\[4\]
+ net126 _1029_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__mux4_1
XANTENNA__5355__S1 _1706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6014_ _2717_ _2752_ _1146_ VGND VGND VPWR VPWR _2753_ sky130_fd_sc_hd__mux2_1
XANTENNA__5680__A1 _1148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8544__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5107__S1 _1708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7965_ net878 _3450_ _3915_ VGND VGND VPWR VPWR _3949_ sky130_fd_sc_hd__mux2_1
XANTENNA__5432__A1 _1686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6916_ _3377_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__clkbuf_1
X_7896_ _3912_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6847_ net674 _3089_ _3340_ VGND VGND VPWR VPWR _3341_ sky130_fd_sc_hd__mux2_1
XANTENNA__7185__A1 _3489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9566_ clknet_leaf_72_clk _0726_ VGND VGND VPWR VPWR rf.registers\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6778_ _3303_ VGND VGND VPWR VPWR _3304_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5291__S0 _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8517_ _4241_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5729_ _2480_ _2481_ VGND VGND VPWR VPWR _2482_ sky130_fd_sc_hd__or2b_1
X_9497_ clknet_leaf_20_clk _0657_ VGND VGND VPWR VPWR rf.registers\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8448_ net417 net14 _4205_ VGND VGND VPWR VPWR _4206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8379_ _4168_ VGND VGND VPWR VPWR _4169_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7623__S _3758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold360 rf.registers\[12\]\[3\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold371 rf.registers\[11\]\[27\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold382 rf.registers\[19\]\[27\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 rf.registers\[16\]\[26\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8454__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1060 rf.registers\[26\]\[11\] VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 rf.registers\[26\]\[30\] VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5379__A _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6702__S _3253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6923__A1 _3101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer5 net86 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_141_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5034__S0 _1719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8428__A1 _3504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4458__A _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5337__S1 _1642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8364__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4905__B _1660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6611__A0 _3060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4848__S0 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7750_ _3835_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4962_ _1702_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6701_ _3262_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7681_ net1052 _3506_ _3794_ VGND VGND VPWR VPWR _3799_ sky130_fd_sc_hd__mux2_1
X_4893_ _1647_ _1648_ _1645_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9420_ clknet_leaf_45_clk _0580_ VGND VGND VPWR VPWR rf.registers\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6632_ _3081_ net1011 _3217_ VGND VGND VPWR VPWR _3226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5273__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9351_ clknet_leaf_65_clk _0511_ VGND VGND VPWR VPWR rf.registers\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6563_ _3188_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5514_ _1828_ _2269_ _1728_ VGND VGND VPWR VPWR _2270_ sky130_fd_sc_hd__a21oi_1
X_8302_ _3011_ net922 _4119_ VGND VGND VPWR VPWR _4128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9282_ clknet_leaf_58_clk _0442_ VGND VGND VPWR VPWR rf.registers\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6494_ _3150_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8233_ _4091_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__clkbuf_1
X_5445_ _2197_ _2200_ _1716_ VGND VGND VPWR VPWR _2201_ sky130_fd_sc_hd__mux2_1
XANTENNA__8539__S _4244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7443__S _3664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4689__C1 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5752__A _2503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8419__A1 _3495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8164_ net371 _3444_ _4047_ VGND VGND VPWR VPWR _4055_ sky130_fd_sc_hd__mux2_1
X_5376_ rf.registers\[8\]\[14\] rf.registers\[9\]\[14\] rf.registers\[10\]\[14\] rf.registers\[11\]\[14\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7115_ _3494_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
X_4327_ _1025_ _1070_ _1077_ _1082_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8095_ _4018_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5328__S1 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7046_ _3447_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4861__C1 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8997_ clknet_leaf_61_clk _0157_ VGND VGND VPWR VPWR rf.registers\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_7948_ _3940_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5500__S1 _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7879_ _3137_ net797 _3902_ VGND VGND VPWR VPWR _3904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6522__S _3157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6905__A1 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9549_ clknet_leaf_44_clk _0709_ VGND VGND VPWR VPWR rf.registers\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold190 rf.registers\[6\]\[0\] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5892__B2 _2621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5644__A1 _1842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8184__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7528__S _3711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6432__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5255__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5007__S0 _1676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5230_ _1984_ _1985_ _1901_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__mux2_1
X_5161_ rf.registers\[4\]\[30\] rf.registers\[5\]\[30\] rf.registers\[6\]\[30\] rf.registers\[7\]\[30\]
+ _1881_ _1883_ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5092_ _1846_ _1847_ _1686_ VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8920_ clknet_leaf_12_clk _0080_ VGND VGND VPWR VPWR rf.registers\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8094__S _4011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4916__A _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6607__S _3206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8851_ clknet_leaf_32_clk _0011_ VGND VGND VPWR VPWR rf.registers\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7802_ net206 _3491_ _3855_ VGND VGND VPWR VPWR _3863_ sky130_fd_sc_hd__mux2_1
XANTENNA__5399__B1 _1655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5994_ _1169_ _2124_ _1875_ VGND VGND VPWR VPWR _2734_ sky130_fd_sc_hd__o21a_1
X_8782_ clknet_leaf_29_clk _0966_ VGND VGND VPWR VPWR rf.registers\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4945_ net1 VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__buf_4
X_7733_ _3826_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7664_ net374 _3489_ _3783_ VGND VGND VPWR VPWR _3790_ sky130_fd_sc_hd__mux2_1
X_4876_ _1630_ _1631_ _1178_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9403_ clknet_leaf_36_clk _0563_ VGND VGND VPWR VPWR rf.registers\[24\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6615_ _3194_ VGND VGND VPWR VPWR _3217_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_119_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7595_ _3753_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6546_ net709 _3134_ _3179_ VGND VGND VPWR VPWR _3180_ sky130_fd_sc_hd__mux2_1
X_9334_ clknet_leaf_25_clk _0494_ VGND VGND VPWR VPWR rf.registers\[21\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8269__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9265_ clknet_leaf_41_clk _0425_ VGND VGND VPWR VPWR rf.registers\[23\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6477_ _3140_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7173__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5428_ _2180_ _2181_ _2182_ _2183_ _1712_ _1716_ VGND VGND VPWR VPWR _2184_ sky130_fd_sc_hd__mux4_1
X_8216_ _4082_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__clkbuf_1
X_9196_ clknet_leaf_49_clk _0356_ VGND VGND VPWR VPWR rf.registers\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5359_ rf.registers\[12\]\[15\] rf.registers\[13\]\[15\] rf.registers\[14\]\[15\]
+ rf.registers\[15\]\[15\] _2113_ _2114_ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__mux4_1
X_8147_ net1044 _3495_ _4036_ VGND VGND VPWR VPWR _4046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8078_ _4009_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7029_ _3437_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4826__A _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5485__S0 _1734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7348__S _3613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5237__S0 _1896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7083__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7811__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6290__A1 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5476__S0 _1675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7790__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4730_ rf.registers\[4\]\[14\] rf.registers\[5\]\[14\] rf.registers\[6\]\[14\] rf.registers\[7\]\[14\]
+ net1161 _1279_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_140_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5228__S0 _1881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4661_ rf.registers\[24\]\[23\] rf.registers\[25\]\[23\] rf.registers\[26\]\[23\]
+ rf.registers\[27\]\[23\] _1351_ _1352_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6400_ net38 VGND VGND VPWR VPWR _3087_ sky130_fd_sc_hd__clkbuf_2
X_7380_ _3043_ net914 _3639_ VGND VGND VPWR VPWR _3640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4592_ _1171_ _1339_ _1347_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_114_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold904 rf.registers\[0\]\[24\] VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__dlygate4sd3_1
X_6331_ _3040_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold915 rf.registers\[8\]\[15\] VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 rf.registers\[22\]\[27\] VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 rf.registers\[30\]\[2\] VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5506__S _1696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold948 rf.registers\[28\]\[9\] VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__dlygate4sd3_1
X_9050_ clknet_leaf_37_clk _0210_ VGND VGND VPWR VPWR rf.registers\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5305__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold959 rf.registers\[14\]\[17\] VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _2952_ _2986_ _2987_ VGND VGND VPWR VPWR _2988_ sky130_fd_sc_hd__and3_1
XANTENNA__5400__S0 _1702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8001_ _3968_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__clkbuf_1
X_5213_ _1965_ _1968_ _1700_ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__mux2_1
XANTENNA__5856__B2 _2408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6193_ _2254_ _2858_ VGND VGND VPWR VPWR _2922_ sky130_fd_sc_hd__or2_1
X_5144_ rf.registers\[0\]\[31\] rf.registers\[1\]\[31\] rf.registers\[2\]\[31\] rf.registers\[3\]\[31\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__mux4_1
XANTENNA__6337__S _3044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5075_ rf.registers\[8\]\[19\] rf.registers\[9\]\[19\] rf.registers\[10\]\[19\] rf.registers\[11\]\[19\]
+ _1689_ _1693_ VGND VGND VPWR VPWR _1831_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8903_ clknet_leaf_1_clk _0063_ VGND VGND VPWR VPWR rf.registers\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_8834_ clknet_leaf_55_clk _1018_ VGND VGND VPWR VPWR rf.registers\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8552__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8765_ clknet_leaf_15_clk _0949_ VGND VGND VPWR VPWR rf.registers\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7781__A1 _3470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5977_ _2697_ _2717_ _1803_ VGND VGND VPWR VPWR _2718_ sky130_fd_sc_hd__mux2_1
XANTENNA__7168__S _3517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7716_ _3817_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__clkbuf_1
X_4928_ _1645_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__buf_4
X_8696_ clknet_leaf_17_clk _0880_ VGND VGND VPWR VPWR rf.registers\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5219__S0 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7647_ net476 _3472_ _3772_ VGND VGND VPWR VPWR _3781_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4859_ rf.registers\[12\]\[19\] rf.registers\[13\]\[19\] rf.registers\[14\]\[19\]
+ rf.registers\[15\]\[19\] _1173_ _1175_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6800__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7578_ _3744_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9317_ clknet_leaf_57_clk _0477_ VGND VGND VPWR VPWR rf.registers\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6529_ net644 _3118_ _3168_ VGND VGND VPWR VPWR _3171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4320__S _1048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9248_ clknet_leaf_69_clk _0408_ VGND VGND VPWR VPWR rf.registers\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9179_ clknet_leaf_22_clk _0339_ VGND VGND VPWR VPWR rf.registers\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__7631__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5940__A _1480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8462__S _4205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5458__S0 _2051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7806__S _3855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6710__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7107__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7541__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5850__A _2229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4466__A _1221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7460__A0 _3056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8372__S _4155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5900_ _2210_ _2632_ VGND VGND VPWR VPWR _2645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6880_ net513 _3126_ _3351_ VGND VGND VPWR VPWR _3358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5831_ _2578_ VGND VGND VPWR VPWR _2579_ sky130_fd_sc_hd__inv_2
XANTENNA__5297__A _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5762_ _2489_ _2494_ _2505_ _2513_ _2408_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__o32a_2
X_8550_ net608 net22 _4255_ VGND VGND VPWR VPWR _4259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4577__B2 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7501_ _3029_ net807 _3700_ VGND VGND VPWR VPWR _3704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4713_ rf.registers\[24\]\[13\] rf.registers\[25\]\[13\] rf.registers\[26\]\[13\]
+ rf.registers\[27\]\[13\] net126 _1029_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__mux4_1
X_5693_ _1145_ net1169 _2411_ VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__a21oi_1
X_8481_ net370 net21 _4216_ VGND VGND VPWR VPWR _4223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7432_ _3667_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__clkbuf_1
X_4644_ rf.registers\[20\]\[7\] rf.registers\[21\]\[7\] rf.registers\[22\]\[7\] rf.registers\[23\]\[7\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__mux4_1
XANTENNA__6620__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4424__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7363_ _3027_ net1073 _3628_ VGND VGND VPWR VPWR _3631_ sky130_fd_sc_hd__mux2_1
Xhold701 rf.registers\[15\]\[14\] VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ rf.registers\[0\]\[31\] rf.registers\[1\]\[31\] rf.registers\[2\]\[31\] rf.registers\[3\]\[31\]
+ _1324_ _1325_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__mux4_1
Xhold712 rf.registers\[6\]\[16\] VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold723 rf.registers\[23\]\[27\] VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd3_1
X_9102_ clknet_leaf_43_clk _0262_ VGND VGND VPWR VPWR rf.registers\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6314_ net39 VGND VGND VPWR VPWR _3029_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold734 rf.registers\[16\]\[15\] VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
X_7294_ _3027_ net796 _3591_ VGND VGND VPWR VPWR _3594_ sky130_fd_sc_hd__mux2_1
Xhold745 rf.registers\[7\]\[24\] VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 rf.registers\[20\]\[8\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 rf.registers\[30\]\[6\] VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 rf.registers\[8\]\[1\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlygate4sd3_1
X_9033_ clknet_leaf_51_clk _0193_ VGND VGND VPWR VPWR rf.registers\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6245_ _2675_ _2703_ _1803_ VGND VGND VPWR VPWR _2971_ sky130_fd_sc_hd__mux2_1
Xhold789 rf.registers\[4\]\[2\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6176_ _2904_ _2905_ VGND VGND VPWR VPWR _2906_ sky130_fd_sc_hd__xnor2_1
X_5127_ _1723_ VGND VGND VPWR VPWR _1883_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5058_ _1812_ _1813_ _1713_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4360__S0 _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8817_ clknet_leaf_43_clk _1001_ VGND VGND VPWR VPWR rf.registers\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_140_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8748_ clknet_leaf_63_clk _0932_ VGND VGND VPWR VPWR rf.registers\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5000__A _1668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4663__S1 _1352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8679_ clknet_leaf_66_clk _0863_ VGND VGND VPWR VPWR rf.registers\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8311__A _4132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5654__B net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5146__S _1901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7361__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6493__A1 _3013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4286__A _1041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold61 rf.registers\[1\]\[9\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 rf.registers\[1\]\[13\] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 rf.registers\[1\]\[26\] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 rf.registers\[0\]\[9\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8192__S _4061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5845__A _1111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4406__S1 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_3 _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4360_ _1112_ _1113_ _1114_ _1115_ _1047_ _1050_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_78_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4291_ net6 VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5580__A _1060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6030_ _1634_ _2767_ VGND VGND VPWR VPWR _2768_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_91_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6236__A1 _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6236__B2 _1127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7981_ _3103_ net982 _3952_ VGND VGND VPWR VPWR _3958_ sky130_fd_sc_hd__mux2_1
Xrebuffer15 _1237_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_109_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer37 net118 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlymetal6s2s_1
X_6932_ _3385_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4924__A _1679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer48 _1217_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
X_6863_ net240 _3109_ _3340_ VGND VGND VPWR VPWR _3349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8602_ clknet_leaf_35_clk _0786_ VGND VGND VPWR VPWR rf.registers\[22\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5814_ _2539_ _2543_ _2562_ VGND VGND VPWR VPWR _2563_ sky130_fd_sc_hd__o21ai_1
X_9582_ clknet_leaf_28_clk _0742_ VGND VGND VPWR VPWR rf.registers\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6794_ _3312_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4645__S1 _1105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8533_ net288 net45 _4244_ VGND VGND VPWR VPWR _4250_ sky130_fd_sc_hd__mux2_1
X_5745_ _2327_ _1169_ _1661_ VGND VGND VPWR VPWR _2497_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5755__A _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8464_ net212 net44 _4205_ VGND VGND VPWR VPWR _4214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5676_ _2428_ _2429_ VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__nor2_1
XANTENNA__5474__B _2229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7415_ _3079_ net1015 _3650_ VGND VGND VPWR VPWR _3658_ sky130_fd_sc_hd__mux2_1
X_4627_ _1254_ _1382_ _1239_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__o21ai_1
X_8395_ _4177_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7970__A _3951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5070__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold520 rf.registers\[11\]\[30\] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold531 rf.registers\[22\]\[28\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _1214_ _1313_ _1239_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__o21ai_1
X_7346_ _3079_ net517 _3613_ VGND VGND VPWR VPWR _3621_ sky130_fd_sc_hd__mux2_1
Xhold542 rf.registers\[24\]\[12\] VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold553 rf.registers\[29\]\[20\] VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 rf.registers\[19\]\[20\] VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__8277__S _4108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold575 rf.registers\[11\]\[24\] VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlygate4sd3_1
X_7277_ _3584_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
X_4489_ _1243_ _1244_ _1211_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__mux2_1
Xhold586 rf.registers\[12\]\[21\] VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7181__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold597 rf.registers\[21\]\[28\] VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9016_ clknet_leaf_12_clk _0176_ VGND VGND VPWR VPWR rf.registers\[31\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6228_ _2953_ _2954_ VGND VGND VPWR VPWR _2955_ sky130_fd_sc_hd__or2_4
XFILLER_0_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6159_ _2015_ _2889_ VGND VGND VPWR VPWR _2890_ sky130_fd_sc_hd__nand2_1
XANTENNA__4581__S0 _1267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__9315__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6525__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5306__A1_N _1729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clone25_A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8152__A1 _3500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5061__S1 _1707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5910__B1 _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput51 net51 VGND VGND VPWR VPWR alu_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__6466__A1 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput62 net62 VGND VGND VPWR VPWR alu_out[21] sky130_fd_sc_hd__buf_2
Xoutput73 net73 VGND VGND VPWR VPWR alu_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_128_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4572__S0 _1324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6218__A1 _2255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6218__B2 _2337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6435__S _3093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4324__S0 _1042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__7120__A _3455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4875__S1 _1175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__8832__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7266__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5575__A _1669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5530_ _1670_ _2277_ _2281_ _2285_ VGND VGND VPWR VPWR _2286_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5461_ rf.registers\[28\]\[8\] rf.registers\[29\]\[8\] rf.registers\[30\]\[8\] rf.registers\[31\]\[8\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5052__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4412_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__buf_2
X_7200_ net556 _3504_ _3539_ VGND VGND VPWR VPWR _3543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8180_ net408 _3460_ _4061_ VGND VGND VPWR VPWR _4064_ sky130_fd_sc_hd__mux2_1
X_5392_ rf.registers\[28\]\[13\] rf.registers\[29\]\[13\] rf.registers\[30\]\[13\]
+ rf.registers\[31\]\[13\] _1673_ _1690_ VGND VGND VPWR VPWR _2148_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4343_ rf.registers\[8\]\[3\] rf.registers\[9\]\[3\] rf.registers\[10\]\[3\] rf.registers\[11\]\[3\]
+ net103 _1044_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7131_ _3505_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4919__A _1674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6457__A1 _3126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7062_ net561 _3458_ _3456_ VGND VGND VPWR VPWR _3459_ sky130_fd_sc_hd__mux2_1
XANTENNA__9338__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4274_ rf.registers\[20\]\[4\] rf.registers\[21\]\[4\] rf.registers\[22\]\[4\] rf.registers\[23\]\[4\]
+ _1027_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6013_ _2341_ _2401_ VGND VGND VPWR VPWR _2752_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4654__A _1071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5968__B1 _2411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
X_7964_ _3948_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6915_ net549 _3089_ _3376_ VGND VGND VPWR VPWR _3377_ sky130_fd_sc_hd__mux2_1
X_7895_ _3013_ net1063 _3902_ VGND VGND VPWR VPWR _3912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8560__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6846_ _3339_ VGND VGND VPWR VPWR _3340_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_wire82_A _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9565_ clknet_leaf_14_clk _0725_ VGND VGND VPWR VPWR rf.registers\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6777_ _3005_ _3302_ VGND VGND VPWR VPWR _3303_ sky130_fd_sc_hd__nor2_4
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8516_ net686 net25 _3007_ VGND VGND VPWR VPWR _4241_ sky130_fd_sc_hd__mux2_1
XANTENNA__5291__S1 _1691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5728_ _2062_ _2479_ VGND VGND VPWR VPWR _2481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9496_ clknet_leaf_27_clk _0656_ VGND VGND VPWR VPWR rf.registers\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8447_ _4204_ VGND VGND VPWR VPWR _4205_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5659_ _2097_ _2410_ _2412_ VGND VGND VPWR VPWR _2414_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7893__A0 _3011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8378_ _3155_ _3192_ VGND VGND VPWR VPWR _4168_ sky130_fd_sc_hd__nor2b_4
Xhold350 rf.registers\[20\]\[3\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold361 rf.registers\[0\]\[14\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
X_7329_ _3062_ net1110 _3602_ VGND VGND VPWR VPWR _3612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold372 rf.registers\[7\]\[1\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6448__A1 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold383 rf.registers\[18\]\[20\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 rf.registers\[2\]\[8\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1050 rf.registers\[25\]\[16\] VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 rf.registers\[24\]\[11\] VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 rf.registers\[21\]\[23\] VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4306__S0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7086__S _3456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer6 _2657_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5034__S1 _1722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5842__B _2040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4739__A _1464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6439__A1 _3113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output63_A net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4545__S0 _1262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6165__S _2327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4474__A _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4848__S1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4961_ _1716_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__buf_4
XANTENNA__8380__S _4169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6700_ net851 _3011_ _3253_ VGND VGND VPWR VPWR _3262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7680_ _3798_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8364__A1 _3508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4892_ rf.registers\[24\]\[0\] rf.registers\[25\]\[0\] rf.registers\[26\]\[0\] rf.registers\[27\]\[0\]
+ net1 net2 VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6631_ _3225_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5509__S _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5273__S1 _1919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9350_ clknet_leaf_0_clk _0510_ VGND VGND VPWR VPWR rf.registers\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6562_ net959 _3011_ _3179_ VGND VGND VPWR VPWR _3188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__8116__A1 _3464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8301_ _4127_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5513_ _2267_ _2268_ _1738_ VGND VGND VPWR VPWR _2269_ sky130_fd_sc_hd__mux2_1
X_9281_ clknet_leaf_56_clk _0441_ VGND VGND VPWR VPWR rf.registers\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6493_ net645 _3013_ _3135_ VGND VGND VPWR VPWR _3150_ sky130_fd_sc_hd__mux2_1
XANTENNA__7724__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8232_ net984 _3444_ _4083_ VGND VGND VPWR VPWR _4091_ sky130_fd_sc_hd__mux2_1
X_5444_ _2198_ _2199_ _2044_ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
X_8163_ _4054_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__clkbuf_1
X_5375_ _2127_ _2130_ _1696_ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7025__A _3412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7114_ net391 _3493_ _3477_ VGND VGND VPWR VPWR _3494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4326_ _1078_ _1081_ _1057_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__a21oi_1
X_8094_ net628 _3442_ _4011_ VGND VGND VPWR VPWR _4018_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_26_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7045_ net858 _3446_ _3435_ VGND VGND VPWR VPWR _3447_ sky130_fd_sc_hd__mux2_1
XANTENNA__4536__S0 _1291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8996_ clknet_leaf_62_clk _0156_ VGND VGND VPWR VPWR rf.registers\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__5405__A2 _2160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7947_ net467 _3500_ _3938_ VGND VGND VPWR VPWR _3940_ sky130_fd_sc_hd__mux2_1
XANTENNA__4613__B1 _1239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__8290__S _4119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7878_ _3903_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_35_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6829_ net936 _3143_ _3326_ VGND VGND VPWR VPWR _3331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9548_ clknet_leaf_45_clk _0708_ VGND VGND VPWR VPWR rf.registers\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6104__A _1754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9479_ clknet_leaf_68_clk _0639_ VGND VGND VPWR VPWR rf.registers\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__6669__A1 _3120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5341__A1 _1640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4775__S0 _1290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold180 rf.registers\[31\]\[23\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold191 rf.registers\[8\]\[10\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4527__S0 net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7809__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5255__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4368__C1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5007__S1 _1681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4766__S0 _1149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5883__A2 _2591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5160_ _1773_ _1915_ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__nor2_1
XANTENNA__4518__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5091_ rf.registers\[24\]\[17\] rf.registers\[25\]\[17\] rf.registers\[26\]\[17\]
+ rf.registers\[27\]\[17\] _1689_ _1693_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__mux4_1
XANTENNA__5191__S0 _1882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4408__S _1035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8850_ clknet_leaf_25_clk _0010_ VGND VGND VPWR VPWR rf.registers\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_7801_ _3862_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5399__A1 _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8781_ clknet_leaf_44_clk _0965_ VGND VGND VPWR VPWR rf.registers\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5993_ _2327_ _2675_ _2732_ VGND VGND VPWR VPWR _2733_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7732_ _3056_ net441 _3819_ VGND VGND VPWR VPWR _3826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4944_ _1699_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7663_ _3789_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4875_ rf.registers\[0\]\[18\] rf.registers\[1\]\[18\] rf.registers\[2\]\[18\] rf.registers\[3\]\[18\]
+ net132 _1175_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6899__A1 _3145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9402_ clknet_leaf_37_clk _0562_ VGND VGND VPWR VPWR rf.registers\[24\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6614_ _3216_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_119_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7594_ _3054_ net1095 _3747_ VGND VGND VPWR VPWR _3753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9333_ clknet_leaf_31_clk _0493_ VGND VGND VPWR VPWR rf.registers\[21\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6545_ _3156_ VGND VGND VPWR VPWR _3179_ sky130_fd_sc_hd__buf_4
XANTENNA__7454__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9264_ clknet_leaf_13_clk _0424_ VGND VGND VPWR VPWR rf.registers\[23\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6476_ net332 _3139_ _3135_ VGND VGND VPWR VPWR _3140_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8215_ net944 _3495_ _4072_ VGND VGND VPWR VPWR _4082_ sky130_fd_sc_hd__mux2_1
X_5427_ rf.registers\[20\]\[11\] rf.registers\[21\]\[11\] rf.registers\[22\]\[11\]
+ rf.registers\[23\]\[11\] _1675_ _1692_ VGND VGND VPWR VPWR _2183_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5323__B2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4757__S0 _1026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9195_ clknet_leaf_2_clk _0355_ VGND VGND VPWR VPWR rf.registers\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8146_ _4045_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__clkbuf_1
X_5358_ _2052_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8273__A0 _3122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4309_ A2[0] VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__buf_12
XANTENNA__6594__A _3194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8077_ net1128 _3493_ _4000_ VGND VGND VPWR VPWR _4009_ sky130_fd_sc_hd__mux2_1
X_5289_ _2042_ _2043_ _2044_ VGND VGND VPWR VPWR _2045_ sky130_fd_sc_hd__mux2_1
XANTENNA__6823__A1 _3137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7028_ net457 _3137_ _3435_ VGND VGND VPWR VPWR _3437_ sky130_fd_sc_hd__mux2_1
XANTENNA__5182__S0 _1767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8979_ clknet_leaf_35_clk _0139_ VGND VGND VPWR VPWR rf.registers\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5485__S1 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6533__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5237__S1 _1898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4988__S _1697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__8500__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4748__S0 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6275__C1 _1087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7539__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5476__S1 _1692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5228__S1 _1883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4660_ _1399_ _1415_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__nand2_4
XFILLER_0_83_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4591_ _1341_ _1343_ _1346_ _1187_ _1215_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__o221a_4
XANTENNA__7274__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5583__A _1167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6330_ _3039_ net587 _3023_ VGND VGND VPWR VPWR _3040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold905 rf.registers\[15\]\[7\] VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold916 rf.registers\[27\]\[14\] VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold927 rf.registers\[5\]\[7\] VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 rf.registers\[26\]\[5\] VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5305__A1 _1699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold949 rf.registers\[14\]\[3\] VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6261_ _2934_ _2940_ _2951_ _2932_ VGND VGND VPWR VPWR _2987_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8000_ _3122_ net1092 _3963_ VGND VGND VPWR VPWR _3968_ sky130_fd_sc_hd__mux2_1
XANTENNA__5400__S1 _1678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5212_ _1966_ _1967_ _1745_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6192_ _2918_ _2920_ VGND VGND VPWR VPWR _2921_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6618__S _3217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5143_ rf.registers\[4\]\[31\] rf.registers\[5\]\[31\] rf.registers\[6\]\[31\] rf.registers\[7\]\[31\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__mux4_1
X_5074_ rf.registers\[12\]\[19\] rf.registers\[13\]\[19\] rf.registers\[14\]\[19\]
+ rf.registers\[15\]\[19\] _1689_ _1693_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__mux4_1
XANTENNA__5164__S0 _1918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4816__B1 _1567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8902_ clknet_leaf_1_clk _0062_ VGND VGND VPWR VPWR rf.registers\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__8558__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8833_ clknet_leaf_53_clk _1017_ VGND VGND VPWR VPWR rf.registers\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5758__A _2305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8764_ clknet_leaf_16_clk _0948_ VGND VGND VPWR VPWR rf.registers\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_5976_ _2344_ _2342_ VGND VGND VPWR VPWR _2717_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_23_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7715_ _3039_ net881 _3808_ VGND VGND VPWR VPWR _3817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4927_ rf.registers\[16\]\[23\] rf.registers\[17\]\[23\] rf.registers\[18\]\[23\]
+ rf.registers\[19\]\[23\] _1676_ _1681_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__mux4_1
X_8695_ clknet_leaf_23_clk _0879_ VGND VGND VPWR VPWR rf.registers\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5219__S1 _1897_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7646_ _3780_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4858_ rf.registers\[8\]\[19\] rf.registers\[9\]\[19\] rf.registers\[10\]\[19\] rf.registers\[11\]\[19\]
+ _1173_ _1175_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6741__A0 _3054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7577_ _3037_ net784 _3736_ VGND VGND VPWR VPWR _3744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4789_ _1543_ _1544_ _1034_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9316_ clknet_leaf_52_clk _0476_ VGND VGND VPWR VPWR rf.registers\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6528_ _3170_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__clkbuf_1
X_9247_ clknet_leaf_73_clk _0407_ VGND VGND VPWR VPWR rf.registers\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6459_ net22 VGND VGND VPWR VPWR _3128_ sky130_fd_sc_hd__buf_2
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9178_ clknet_leaf_17_clk _0338_ VGND VGND VPWR VPWR rf.registers\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__8246__A0 _3095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8129_ net500 _3476_ _4036_ VGND VGND VPWR VPWR _4037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7359__S _3628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5458__S1 _2053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4969__S0 _1720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7123__A net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7212__A1 _3448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5830_ _2577_ _2498_ _1803_ VGND VGND VPWR VPWR _2578_ sky130_fd_sc_hd__mux2_1
XANTENNA__4482__A _1217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5761_ _2511_ _2512_ VGND VGND VPWR VPWR _2513_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7500_ _3703_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4712_ rf.registers\[28\]\[13\] rf.registers\[29\]\[13\] rf.registers\[30\]\[13\]
+ rf.registers\[31\]\[13\] net126 _1029_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6901__S _3362_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8480_ _4222_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__clkbuf_1
X_5692_ _1666_ _2445_ VGND VGND VPWR VPWR _2446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7431_ _3027_ net973 _3664_ VGND VGND VPWR VPWR _3667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4643_ _1025_ _1390_ _1398_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7362_ _3630_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6202__A _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4574_ rf.registers\[4\]\[31\] rf.registers\[5\]\[31\] rf.registers\[6\]\[31\] rf.registers\[7\]\[31\]
+ _1324_ _1325_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__mux4_1
Xhold702 rf.registers\[28\]\[7\] VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 rf.registers\[31\]\[8\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd3_1
X_9101_ clknet_leaf_50_clk _0261_ VGND VGND VPWR VPWR rf.registers\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold724 rf.registers\[31\]\[3\] VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ _3028_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold735 rf.registers\[24\]\[20\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 rf.registers\[2\]\[7\] VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd3_1
X_7293_ _3593_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7732__S _3819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold757 rf.registers\[6\]\[23\] VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 rf.registers\[24\]\[0\] VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__dlygate4sd3_1
X_9032_ clknet_leaf_46_clk _0192_ VGND VGND VPWR VPWR rf.registers\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold779 rf.registers\[27\]\[6\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ _2672_ _2674_ _1803_ VGND VGND VPWR VPWR _2970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6175_ _2887_ _2890_ _2892_ VGND VGND VPWR VPWR _2905_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5126_ _1881_ VGND VGND VPWR VPWR _1882_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_127_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5057_ rf.registers\[12\]\[18\] rf.registers\[13\]\[18\] rf.registers\[14\]\[18\]
+ rf.registers\[15\]\[18\] _1689_ _1693_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__mux4_1
XANTENNA__4360__S1 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7179__S _3528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_8816_ clknet_leaf_12_clk _1000_ VGND VGND VPWR VPWR rf.registers\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8747_ clknet_leaf_4_clk _0931_ VGND VGND VPWR VPWR rf.registers\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5959_ _2335_ _2701_ VGND VGND VPWR VPWR _2702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7907__S _3916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8678_ clknet_leaf_1_clk _0862_ VGND VGND VPWR VPWR rf.registers\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5935__B net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7629_ _3005_ _3153_ VGND VGND VPWR VPWR _3771_ sky130_fd_sc_hd__nor2_4
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6112__A _2102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5376__S0 _2113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8039__A _3988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold62 rf.registers\[1\]\[25\] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold73 rf.registers\[18\]\[12\] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8473__S _4216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold84 rf.registers\[24\]\[13\] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 rf.registers\[6\]\[10\] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5453__B1 _1728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7817__S _3866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__8611__CLK clknet_leaf_68_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _1717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4290_ _1040_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5580__B _1085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_6_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7980_ _3957_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5800__S _2501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer16 net97 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_109_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6931_ net1047 _3109_ _3376_ VGND VGND VPWR VPWR _3385_ sky130_fd_sc_hd__mux2_1
Xrebuffer38 _2661_ VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer49 _2535_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6862_ _3348_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8601_ clknet_leaf_19_clk _0785_ VGND VGND VPWR VPWR rf.registers\[22\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5813_ _2271_ _2538_ VGND VGND VPWR VPWR _2562_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9581_ clknet_leaf_44_clk _0741_ VGND VGND VPWR VPWR rf.registers\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6793_ net813 _3107_ _3304_ VGND VGND VPWR VPWR _3312_ sky130_fd_sc_hd__mux2_1
XANTENNA__9267__CLK clknet_leaf_35_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8532_ _4249_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4940__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5744_ _2495_ VGND VGND VPWR VPWR _2496_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_98_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8463_ _4213_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__clkbuf_1
X_5675_ _1800_ _2247_ VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7414_ _3657_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4707__C1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4626_ _1380_ _1381_ _1190_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__mux2_1
X_8394_ net353 _3470_ _4169_ VGND VGND VPWR VPWR _4177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold510 rf.registers\[6\]\[29\] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7345_ _3620_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6867__A _3339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold521 rf.registers\[30\]\[31\] VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8558__S _4255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4557_ _1311_ _1312_ _1199_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__mux2_1
Xhold532 rf.registers\[21\]\[13\] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7462__S _3675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold543 rf.registers\[29\]\[19\] VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 rf.registers\[28\]\[11\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold565 rf.registers\[11\]\[22\] VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__dlygate4sd3_1
X_7276_ _3077_ net630 _3577_ VGND VGND VPWR VPWR _3584_ sky130_fd_sc_hd__mux2_1
Xhold576 rf.registers\[0\]\[17\] VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ rf.registers\[24\]\[20\] rf.registers\[25\]\[20\] rf.registers\[26\]\[20\]
+ rf.registers\[27\]\[20\] _1207_ _1208_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__mux4_1
Xhold587 rf.registers\[11\]\[7\] VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 rf.registers\[22\]\[0\] VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__dlygate4sd3_1
X_9015_ clknet_leaf_33_clk _0175_ VGND VGND VPWR VPWR rf.registers\[31\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6227_ _2940_ _2934_ _2932_ VGND VGND VPWR VPWR _2954_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_129_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _1370_ _2888_ VGND VGND VPWR VPWR _2889_ sky130_fd_sc_hd__xor2_1
XANTENNA__4581__S1 _1268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7698__A _3807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5109_ _1861_ _1862_ _1863_ _1864_ _1713_ _1717_ VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_142_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6806__S _3315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6089_ _2756_ _2751_ _2426_ VGND VGND VPWR VPWR _2824_ sky130_fd_sc_hd__mux2_1
XANTENNA__5710__S _2178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5011__A _1704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7637__S _3772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6541__S _3168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4410__A1 _1057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clone18_A _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4996__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput52 net52 VGND VGND VPWR VPWR alu_out[12] sky130_fd_sc_hd__buf_6
Xoutput63 net63 VGND VGND VPWR VPWR alu_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__4297__A _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput74 net74 VGND VGND VPWR VPWR alu_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_101_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4572__S1 _1325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6716__S _3267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5521__S0 _1711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4324__S1 _1044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7547__S _3722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6451__S _3114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5575__B _1660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5460_ _2214_ _2215_ _1685_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4411_ net1170 VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__buf_2
XFILLER_0_112_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5391_ _2145_ _2146_ _1684_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7282__S _3577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7130_ net329 _3504_ _3498_ VGND VGND VPWR VPWR _3505_ sky130_fd_sc_hd__mux2_1
X_4342_ _1038_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__7654__A1 _3479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7061_ net25 VGND VGND VPWR VPWR _3458_ sky130_fd_sc_hd__buf_2
X_4273_ _1028_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__buf_4
X_6012_ _2649_ _2697_ _2327_ VGND VGND VPWR VPWR _2751_ sky130_fd_sc_hd__mux2_1
.ends

