VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 434.795 BY 445.515 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END A1[4]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.368000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.886500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END A2[4]
  PIN A3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END A3[4]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 10.640 39.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.020 10.640 64.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.020 10.640 89.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.020 10.640 114.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.020 10.640 139.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 163.020 10.640 164.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 10.640 189.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.020 10.640 214.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 238.020 10.640 239.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.020 10.640 264.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.020 10.640 289.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 313.020 10.640 314.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.020 10.640 339.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 363.020 10.640 364.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 388.020 10.640 389.620 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.020 10.640 414.620 432.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.380 429.420 19.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.380 429.420 44.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.380 429.420 69.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 93.380 429.420 94.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 118.380 429.420 119.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 143.380 429.420 144.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 168.380 429.420 169.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 193.380 429.420 194.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 218.380 429.420 219.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 243.380 429.420 244.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 268.380 429.420 269.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 293.380 429.420 294.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 318.380 429.420 319.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 343.380 429.420 344.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 368.380 429.420 369.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 393.380 429.420 394.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 418.380 429.420 419.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.720 10.640 61.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.720 10.640 86.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 109.720 10.640 111.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.720 10.640 136.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.720 10.640 161.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 10.640 186.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.720 10.640 211.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.720 10.640 236.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 259.720 10.640 261.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.720 10.640 286.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 309.720 10.640 311.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.720 10.640 336.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 359.720 10.640 361.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.720 10.640 386.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 409.720 10.640 411.320 432.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 429.420 16.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.080 429.420 41.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 65.080 429.420 66.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 90.080 429.420 91.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 115.080 429.420 116.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 140.080 429.420 141.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 165.080 429.420 166.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 190.080 429.420 191.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 215.080 429.420 216.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 240.080 429.420 241.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 265.080 429.420 266.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 290.080 429.420 291.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 315.080 429.420 316.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 340.080 429.420 341.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 365.080 429.420 366.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 390.080 429.420 391.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 415.080 429.420 416.680 ;
    END
  END VPWR
  PIN WD3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END WD3[0]
  PIN WD3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END WD3[10]
  PIN WD3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END WD3[11]
  PIN WD3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END WD3[12]
  PIN WD3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END WD3[13]
  PIN WD3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END WD3[14]
  PIN WD3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END WD3[15]
  PIN WD3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END WD3[16]
  PIN WD3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END WD3[17]
  PIN WD3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END WD3[18]
  PIN WD3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END WD3[19]
  PIN WD3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END WD3[1]
  PIN WD3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END WD3[20]
  PIN WD3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END WD3[21]
  PIN WD3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END WD3[22]
  PIN WD3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END WD3[23]
  PIN WD3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END WD3[24]
  PIN WD3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END WD3[25]
  PIN WD3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END WD3[26]
  PIN WD3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END WD3[27]
  PIN WD3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END WD3[28]
  PIN WD3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END WD3[29]
  PIN WD3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END WD3[2]
  PIN WD3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END WD3[30]
  PIN WD3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END WD3[31]
  PIN WD3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END WD3[3]
  PIN WD3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END WD3[4]
  PIN WD3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END WD3[5]
  PIN WD3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END WD3[6]
  PIN WD3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END WD3[7]
  PIN WD3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END WD3[8]
  PIN WD3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END WD3[9]
  PIN WE3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END WE3
  PIN alu_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 10.920 434.795 11.520 ;
    END
  END alu_out[0]
  PIN alu_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 146.920 434.795 147.520 ;
    END
  END alu_out[10]
  PIN alu_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 160.520 434.795 161.120 ;
    END
  END alu_out[11]
  PIN alu_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 174.120 434.795 174.720 ;
    END
  END alu_out[12]
  PIN alu_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 187.720 434.795 188.320 ;
    END
  END alu_out[13]
  PIN alu_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 201.320 434.795 201.920 ;
    END
  END alu_out[14]
  PIN alu_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 214.920 434.795 215.520 ;
    END
  END alu_out[15]
  PIN alu_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 430.795 228.520 434.795 229.120 ;
    END
  END alu_out[16]
  PIN alu_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 242.120 434.795 242.720 ;
    END
  END alu_out[17]
  PIN alu_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 430.795 255.720 434.795 256.320 ;
    END
  END alu_out[18]
  PIN alu_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 269.320 434.795 269.920 ;
    END
  END alu_out[19]
  PIN alu_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 24.520 434.795 25.120 ;
    END
  END alu_out[1]
  PIN alu_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 282.920 434.795 283.520 ;
    END
  END alu_out[20]
  PIN alu_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 296.520 434.795 297.120 ;
    END
  END alu_out[21]
  PIN alu_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 310.120 434.795 310.720 ;
    END
  END alu_out[22]
  PIN alu_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 323.720 434.795 324.320 ;
    END
  END alu_out[23]
  PIN alu_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 337.320 434.795 337.920 ;
    END
  END alu_out[24]
  PIN alu_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 350.920 434.795 351.520 ;
    END
  END alu_out[25]
  PIN alu_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 364.520 434.795 365.120 ;
    END
  END alu_out[26]
  PIN alu_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 378.120 434.795 378.720 ;
    END
  END alu_out[27]
  PIN alu_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 391.720 434.795 392.320 ;
    END
  END alu_out[28]
  PIN alu_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 405.320 434.795 405.920 ;
    END
  END alu_out[29]
  PIN alu_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 430.795 38.120 434.795 38.720 ;
    END
  END alu_out[2]
  PIN alu_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 430.795 418.920 434.795 419.520 ;
    END
  END alu_out[30]
  PIN alu_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 432.520 434.795 433.120 ;
    END
  END alu_out[31]
  PIN alu_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 51.720 434.795 52.320 ;
    END
  END alu_out[3]
  PIN alu_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 65.320 434.795 65.920 ;
    END
  END alu_out[4]
  PIN alu_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 78.920 434.795 79.520 ;
    END
  END alu_out[5]
  PIN alu_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 430.795 92.520 434.795 93.120 ;
    END
  END alu_out[6]
  PIN alu_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 106.120 434.795 106.720 ;
    END
  END alu_out[7]
  PIN alu_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 119.720 434.795 120.320 ;
    END
  END alu_out[8]
  PIN alu_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.795 133.320 434.795 133.920 ;
    END
  END alu_out[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END clk
  PIN opcode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END opcode[0]
  PIN opcode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END opcode[1]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 429.370 432.670 ;
      LAYER li1 ;
        RECT 5.520 10.795 429.180 432.565 ;
      LAYER met1 ;
        RECT 0.070 8.880 429.180 438.220 ;
      LAYER met2 ;
        RECT 0.090 8.850 427.250 438.250 ;
      LAYER met3 ;
        RECT 0.065 433.520 430.795 436.385 ;
        RECT 0.065 432.120 430.395 433.520 ;
        RECT 0.065 426.720 430.795 432.120 ;
        RECT 4.400 425.320 430.795 426.720 ;
        RECT 0.065 419.920 430.795 425.320 ;
        RECT 0.065 418.560 430.395 419.920 ;
        RECT 4.400 418.520 430.395 418.560 ;
        RECT 4.400 417.160 430.795 418.520 ;
        RECT 0.065 410.400 430.795 417.160 ;
        RECT 4.400 409.000 430.795 410.400 ;
        RECT 0.065 406.320 430.795 409.000 ;
        RECT 0.065 404.920 430.395 406.320 ;
        RECT 0.065 402.240 430.795 404.920 ;
        RECT 4.400 400.840 430.795 402.240 ;
        RECT 0.065 394.080 430.795 400.840 ;
        RECT 4.400 392.720 430.795 394.080 ;
        RECT 4.400 392.680 430.395 392.720 ;
        RECT 0.065 391.320 430.395 392.680 ;
        RECT 0.065 385.920 430.795 391.320 ;
        RECT 4.400 384.520 430.795 385.920 ;
        RECT 0.065 379.120 430.795 384.520 ;
        RECT 0.065 377.760 430.395 379.120 ;
        RECT 4.400 377.720 430.395 377.760 ;
        RECT 4.400 376.360 430.795 377.720 ;
        RECT 0.065 369.600 430.795 376.360 ;
        RECT 4.400 368.200 430.795 369.600 ;
        RECT 0.065 365.520 430.795 368.200 ;
        RECT 0.065 364.120 430.395 365.520 ;
        RECT 0.065 361.440 430.795 364.120 ;
        RECT 4.400 360.040 430.795 361.440 ;
        RECT 0.065 353.280 430.795 360.040 ;
        RECT 4.400 351.920 430.795 353.280 ;
        RECT 4.400 351.880 430.395 351.920 ;
        RECT 0.065 350.520 430.395 351.880 ;
        RECT 0.065 345.120 430.795 350.520 ;
        RECT 4.400 343.720 430.795 345.120 ;
        RECT 0.065 338.320 430.795 343.720 ;
        RECT 0.065 336.960 430.395 338.320 ;
        RECT 4.400 336.920 430.395 336.960 ;
        RECT 4.400 335.560 430.795 336.920 ;
        RECT 0.065 328.800 430.795 335.560 ;
        RECT 4.400 327.400 430.795 328.800 ;
        RECT 0.065 324.720 430.795 327.400 ;
        RECT 0.065 323.320 430.395 324.720 ;
        RECT 0.065 320.640 430.795 323.320 ;
        RECT 4.400 319.240 430.795 320.640 ;
        RECT 0.065 312.480 430.795 319.240 ;
        RECT 4.400 311.120 430.795 312.480 ;
        RECT 4.400 311.080 430.395 311.120 ;
        RECT 0.065 309.720 430.395 311.080 ;
        RECT 0.065 304.320 430.795 309.720 ;
        RECT 4.400 302.920 430.795 304.320 ;
        RECT 0.065 297.520 430.795 302.920 ;
        RECT 0.065 296.160 430.395 297.520 ;
        RECT 4.400 296.120 430.395 296.160 ;
        RECT 4.400 294.760 430.795 296.120 ;
        RECT 0.065 288.000 430.795 294.760 ;
        RECT 4.400 286.600 430.795 288.000 ;
        RECT 0.065 283.920 430.795 286.600 ;
        RECT 0.065 282.520 430.395 283.920 ;
        RECT 0.065 279.840 430.795 282.520 ;
        RECT 4.400 278.440 430.795 279.840 ;
        RECT 0.065 271.680 430.795 278.440 ;
        RECT 4.400 270.320 430.795 271.680 ;
        RECT 4.400 270.280 430.395 270.320 ;
        RECT 0.065 268.920 430.395 270.280 ;
        RECT 0.065 263.520 430.795 268.920 ;
        RECT 4.400 262.120 430.795 263.520 ;
        RECT 0.065 256.720 430.795 262.120 ;
        RECT 0.065 255.360 430.395 256.720 ;
        RECT 4.400 255.320 430.395 255.360 ;
        RECT 4.400 253.960 430.795 255.320 ;
        RECT 0.065 247.200 430.795 253.960 ;
        RECT 4.400 245.800 430.795 247.200 ;
        RECT 0.065 243.120 430.795 245.800 ;
        RECT 0.065 241.720 430.395 243.120 ;
        RECT 0.065 239.040 430.795 241.720 ;
        RECT 4.400 237.640 430.795 239.040 ;
        RECT 0.065 230.880 430.795 237.640 ;
        RECT 4.400 229.520 430.795 230.880 ;
        RECT 4.400 229.480 430.395 229.520 ;
        RECT 0.065 228.120 430.395 229.480 ;
        RECT 0.065 222.720 430.795 228.120 ;
        RECT 4.400 221.320 430.795 222.720 ;
        RECT 0.065 215.920 430.795 221.320 ;
        RECT 0.065 214.560 430.395 215.920 ;
        RECT 4.400 214.520 430.395 214.560 ;
        RECT 4.400 213.160 430.795 214.520 ;
        RECT 0.065 206.400 430.795 213.160 ;
        RECT 4.400 205.000 430.795 206.400 ;
        RECT 0.065 202.320 430.795 205.000 ;
        RECT 0.065 200.920 430.395 202.320 ;
        RECT 0.065 198.240 430.795 200.920 ;
        RECT 4.400 196.840 430.795 198.240 ;
        RECT 0.065 190.080 430.795 196.840 ;
        RECT 4.400 188.720 430.795 190.080 ;
        RECT 4.400 188.680 430.395 188.720 ;
        RECT 0.065 187.320 430.395 188.680 ;
        RECT 0.065 181.920 430.795 187.320 ;
        RECT 4.400 180.520 430.795 181.920 ;
        RECT 0.065 175.120 430.795 180.520 ;
        RECT 0.065 173.760 430.395 175.120 ;
        RECT 4.400 173.720 430.395 173.760 ;
        RECT 4.400 172.360 430.795 173.720 ;
        RECT 0.065 165.600 430.795 172.360 ;
        RECT 4.400 164.200 430.795 165.600 ;
        RECT 0.065 161.520 430.795 164.200 ;
        RECT 0.065 160.120 430.395 161.520 ;
        RECT 0.065 157.440 430.795 160.120 ;
        RECT 4.400 156.040 430.795 157.440 ;
        RECT 0.065 149.280 430.795 156.040 ;
        RECT 4.400 147.920 430.795 149.280 ;
        RECT 4.400 147.880 430.395 147.920 ;
        RECT 0.065 146.520 430.395 147.880 ;
        RECT 0.065 141.120 430.795 146.520 ;
        RECT 4.400 139.720 430.795 141.120 ;
        RECT 0.065 134.320 430.795 139.720 ;
        RECT 0.065 132.960 430.395 134.320 ;
        RECT 4.400 132.920 430.395 132.960 ;
        RECT 4.400 131.560 430.795 132.920 ;
        RECT 0.065 124.800 430.795 131.560 ;
        RECT 4.400 123.400 430.795 124.800 ;
        RECT 0.065 120.720 430.795 123.400 ;
        RECT 0.065 119.320 430.395 120.720 ;
        RECT 0.065 116.640 430.795 119.320 ;
        RECT 4.400 115.240 430.795 116.640 ;
        RECT 0.065 108.480 430.795 115.240 ;
        RECT 4.400 107.120 430.795 108.480 ;
        RECT 4.400 107.080 430.395 107.120 ;
        RECT 0.065 105.720 430.395 107.080 ;
        RECT 0.065 100.320 430.795 105.720 ;
        RECT 4.400 98.920 430.795 100.320 ;
        RECT 0.065 93.520 430.795 98.920 ;
        RECT 0.065 92.160 430.395 93.520 ;
        RECT 4.400 92.120 430.395 92.160 ;
        RECT 4.400 90.760 430.795 92.120 ;
        RECT 0.065 84.000 430.795 90.760 ;
        RECT 4.400 82.600 430.795 84.000 ;
        RECT 0.065 79.920 430.795 82.600 ;
        RECT 0.065 78.520 430.395 79.920 ;
        RECT 0.065 75.840 430.795 78.520 ;
        RECT 4.400 74.440 430.795 75.840 ;
        RECT 0.065 67.680 430.795 74.440 ;
        RECT 4.400 66.320 430.795 67.680 ;
        RECT 4.400 66.280 430.395 66.320 ;
        RECT 0.065 64.920 430.395 66.280 ;
        RECT 0.065 59.520 430.795 64.920 ;
        RECT 4.400 58.120 430.795 59.520 ;
        RECT 0.065 52.720 430.795 58.120 ;
        RECT 0.065 51.360 430.395 52.720 ;
        RECT 4.400 51.320 430.395 51.360 ;
        RECT 4.400 49.960 430.795 51.320 ;
        RECT 0.065 43.200 430.795 49.960 ;
        RECT 4.400 41.800 430.795 43.200 ;
        RECT 0.065 39.120 430.795 41.800 ;
        RECT 0.065 37.720 430.395 39.120 ;
        RECT 0.065 35.040 430.795 37.720 ;
        RECT 4.400 33.640 430.795 35.040 ;
        RECT 0.065 26.880 430.795 33.640 ;
        RECT 4.400 25.520 430.795 26.880 ;
        RECT 4.400 25.480 430.395 25.520 ;
        RECT 0.065 24.120 430.395 25.480 ;
        RECT 0.065 18.720 430.795 24.120 ;
        RECT 4.400 17.320 430.795 18.720 ;
        RECT 0.065 11.920 430.795 17.320 ;
        RECT 0.065 10.520 430.395 11.920 ;
        RECT 0.065 9.695 430.795 10.520 ;
      LAYER met4 ;
        RECT 0.790 433.120 333.665 436.385 ;
        RECT 0.790 10.240 9.320 433.120 ;
        RECT 11.720 10.240 12.620 433.120 ;
        RECT 15.020 10.240 34.320 433.120 ;
        RECT 36.720 10.240 37.620 433.120 ;
        RECT 40.020 10.240 59.320 433.120 ;
        RECT 61.720 10.240 62.620 433.120 ;
        RECT 65.020 10.240 84.320 433.120 ;
        RECT 86.720 10.240 87.620 433.120 ;
        RECT 90.020 10.240 109.320 433.120 ;
        RECT 111.720 10.240 112.620 433.120 ;
        RECT 115.020 10.240 134.320 433.120 ;
        RECT 136.720 10.240 137.620 433.120 ;
        RECT 140.020 10.240 159.320 433.120 ;
        RECT 161.720 10.240 162.620 433.120 ;
        RECT 165.020 10.240 184.320 433.120 ;
        RECT 186.720 10.240 187.620 433.120 ;
        RECT 190.020 10.240 209.320 433.120 ;
        RECT 211.720 10.240 212.620 433.120 ;
        RECT 215.020 10.240 234.320 433.120 ;
        RECT 236.720 10.240 237.620 433.120 ;
        RECT 240.020 10.240 259.320 433.120 ;
        RECT 261.720 10.240 262.620 433.120 ;
        RECT 265.020 10.240 284.320 433.120 ;
        RECT 286.720 10.240 287.620 433.120 ;
        RECT 290.020 10.240 309.320 433.120 ;
        RECT 311.720 10.240 312.620 433.120 ;
        RECT 315.020 10.240 333.665 433.120 ;
        RECT 0.790 9.695 333.665 10.240 ;
      LAYER met5 ;
        RECT 0.580 421.580 291.980 427.500 ;
        RECT 0.580 413.480 3.680 421.580 ;
        RECT 0.580 396.580 291.980 413.480 ;
        RECT 0.580 388.480 3.680 396.580 ;
        RECT 0.580 371.580 291.980 388.480 ;
        RECT 0.580 363.480 3.680 371.580 ;
        RECT 0.580 346.580 291.980 363.480 ;
        RECT 0.580 338.480 3.680 346.580 ;
        RECT 0.580 321.580 291.980 338.480 ;
        RECT 0.580 313.480 3.680 321.580 ;
        RECT 0.580 296.580 291.980 313.480 ;
        RECT 0.580 288.480 3.680 296.580 ;
        RECT 0.580 271.580 291.980 288.480 ;
        RECT 0.580 263.480 3.680 271.580 ;
        RECT 0.580 246.580 291.980 263.480 ;
        RECT 0.580 238.480 3.680 246.580 ;
        RECT 0.580 221.580 291.980 238.480 ;
        RECT 0.580 213.480 3.680 221.580 ;
        RECT 0.580 196.580 291.980 213.480 ;
        RECT 0.580 188.480 3.680 196.580 ;
        RECT 0.580 171.580 291.980 188.480 ;
        RECT 0.580 163.480 3.680 171.580 ;
        RECT 0.580 146.580 291.980 163.480 ;
        RECT 0.580 138.480 3.680 146.580 ;
        RECT 0.580 121.580 291.980 138.480 ;
        RECT 0.580 113.480 3.680 121.580 ;
        RECT 0.580 96.580 291.980 113.480 ;
        RECT 0.580 88.480 3.680 96.580 ;
        RECT 0.580 71.580 291.980 88.480 ;
        RECT 0.580 63.480 3.680 71.580 ;
        RECT 0.580 48.500 291.980 63.480 ;
  END
END top
END LIBRARY

