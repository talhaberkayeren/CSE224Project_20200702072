module top (WE3,
    clk,
    A1,
    A2,
    A3,
    WD3,
    alu_out,
    opcode);
 input WE3;
 input clk;
 input [4:0] A1;
 input [4:0] A2;
 input [4:0] A3;
 input [31:0] WD3;
 output [31:0] alu_out;
 input [1:0] opcode;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire \rf.registers[0][0] ;
 wire \rf.registers[0][10] ;
 wire \rf.registers[0][11] ;
 wire \rf.registers[0][12] ;
 wire \rf.registers[0][13] ;
 wire \rf.registers[0][14] ;
 wire \rf.registers[0][15] ;
 wire \rf.registers[0][16] ;
 wire \rf.registers[0][17] ;
 wire \rf.registers[0][18] ;
 wire \rf.registers[0][19] ;
 wire \rf.registers[0][1] ;
 wire \rf.registers[0][20] ;
 wire \rf.registers[0][21] ;
 wire \rf.registers[0][22] ;
 wire \rf.registers[0][23] ;
 wire \rf.registers[0][24] ;
 wire \rf.registers[0][25] ;
 wire \rf.registers[0][26] ;
 wire \rf.registers[0][27] ;
 wire \rf.registers[0][28] ;
 wire \rf.registers[0][29] ;
 wire \rf.registers[0][2] ;
 wire \rf.registers[0][30] ;
 wire \rf.registers[0][31] ;
 wire \rf.registers[0][3] ;
 wire \rf.registers[0][4] ;
 wire \rf.registers[0][5] ;
 wire \rf.registers[0][6] ;
 wire \rf.registers[0][7] ;
 wire \rf.registers[0][8] ;
 wire \rf.registers[0][9] ;
 wire \rf.registers[10][0] ;
 wire \rf.registers[10][10] ;
 wire \rf.registers[10][11] ;
 wire \rf.registers[10][12] ;
 wire \rf.registers[10][13] ;
 wire \rf.registers[10][14] ;
 wire \rf.registers[10][15] ;
 wire \rf.registers[10][16] ;
 wire \rf.registers[10][17] ;
 wire \rf.registers[10][18] ;
 wire \rf.registers[10][19] ;
 wire \rf.registers[10][1] ;
 wire \rf.registers[10][20] ;
 wire \rf.registers[10][21] ;
 wire \rf.registers[10][22] ;
 wire \rf.registers[10][23] ;
 wire \rf.registers[10][24] ;
 wire \rf.registers[10][25] ;
 wire \rf.registers[10][26] ;
 wire \rf.registers[10][27] ;
 wire \rf.registers[10][28] ;
 wire \rf.registers[10][29] ;
 wire \rf.registers[10][2] ;
 wire \rf.registers[10][30] ;
 wire \rf.registers[10][31] ;
 wire \rf.registers[10][3] ;
 wire \rf.registers[10][4] ;
 wire \rf.registers[10][5] ;
 wire \rf.registers[10][6] ;
 wire \rf.registers[10][7] ;
 wire \rf.registers[10][8] ;
 wire \rf.registers[10][9] ;
 wire \rf.registers[11][0] ;
 wire \rf.registers[11][10] ;
 wire \rf.registers[11][11] ;
 wire \rf.registers[11][12] ;
 wire \rf.registers[11][13] ;
 wire \rf.registers[11][14] ;
 wire \rf.registers[11][15] ;
 wire \rf.registers[11][16] ;
 wire \rf.registers[11][17] ;
 wire \rf.registers[11][18] ;
 wire \rf.registers[11][19] ;
 wire \rf.registers[11][1] ;
 wire \rf.registers[11][20] ;
 wire \rf.registers[11][21] ;
 wire \rf.registers[11][22] ;
 wire \rf.registers[11][23] ;
 wire \rf.registers[11][24] ;
 wire \rf.registers[11][25] ;
 wire \rf.registers[11][26] ;
 wire \rf.registers[11][27] ;
 wire \rf.registers[11][28] ;
 wire \rf.registers[11][29] ;
 wire \rf.registers[11][2] ;
 wire \rf.registers[11][30] ;
 wire \rf.registers[11][31] ;
 wire \rf.registers[11][3] ;
 wire \rf.registers[11][4] ;
 wire \rf.registers[11][5] ;
 wire \rf.registers[11][6] ;
 wire \rf.registers[11][7] ;
 wire \rf.registers[11][8] ;
 wire \rf.registers[11][9] ;
 wire \rf.registers[12][0] ;
 wire \rf.registers[12][10] ;
 wire \rf.registers[12][11] ;
 wire \rf.registers[12][12] ;
 wire \rf.registers[12][13] ;
 wire \rf.registers[12][14] ;
 wire \rf.registers[12][15] ;
 wire \rf.registers[12][16] ;
 wire \rf.registers[12][17] ;
 wire \rf.registers[12][18] ;
 wire \rf.registers[12][19] ;
 wire \rf.registers[12][1] ;
 wire \rf.registers[12][20] ;
 wire \rf.registers[12][21] ;
 wire \rf.registers[12][22] ;
 wire \rf.registers[12][23] ;
 wire \rf.registers[12][24] ;
 wire \rf.registers[12][25] ;
 wire \rf.registers[12][26] ;
 wire \rf.registers[12][27] ;
 wire \rf.registers[12][28] ;
 wire \rf.registers[12][29] ;
 wire \rf.registers[12][2] ;
 wire \rf.registers[12][30] ;
 wire \rf.registers[12][31] ;
 wire \rf.registers[12][3] ;
 wire \rf.registers[12][4] ;
 wire \rf.registers[12][5] ;
 wire \rf.registers[12][6] ;
 wire \rf.registers[12][7] ;
 wire \rf.registers[12][8] ;
 wire \rf.registers[12][9] ;
 wire \rf.registers[13][0] ;
 wire \rf.registers[13][10] ;
 wire \rf.registers[13][11] ;
 wire \rf.registers[13][12] ;
 wire \rf.registers[13][13] ;
 wire \rf.registers[13][14] ;
 wire \rf.registers[13][15] ;
 wire \rf.registers[13][16] ;
 wire \rf.registers[13][17] ;
 wire \rf.registers[13][18] ;
 wire \rf.registers[13][19] ;
 wire \rf.registers[13][1] ;
 wire \rf.registers[13][20] ;
 wire \rf.registers[13][21] ;
 wire \rf.registers[13][22] ;
 wire \rf.registers[13][23] ;
 wire \rf.registers[13][24] ;
 wire \rf.registers[13][25] ;
 wire \rf.registers[13][26] ;
 wire \rf.registers[13][27] ;
 wire \rf.registers[13][28] ;
 wire \rf.registers[13][29] ;
 wire \rf.registers[13][2] ;
 wire \rf.registers[13][30] ;
 wire \rf.registers[13][31] ;
 wire \rf.registers[13][3] ;
 wire \rf.registers[13][4] ;
 wire \rf.registers[13][5] ;
 wire \rf.registers[13][6] ;
 wire \rf.registers[13][7] ;
 wire \rf.registers[13][8] ;
 wire \rf.registers[13][9] ;
 wire \rf.registers[14][0] ;
 wire \rf.registers[14][10] ;
 wire \rf.registers[14][11] ;
 wire \rf.registers[14][12] ;
 wire \rf.registers[14][13] ;
 wire \rf.registers[14][14] ;
 wire \rf.registers[14][15] ;
 wire \rf.registers[14][16] ;
 wire \rf.registers[14][17] ;
 wire \rf.registers[14][18] ;
 wire \rf.registers[14][19] ;
 wire \rf.registers[14][1] ;
 wire \rf.registers[14][20] ;
 wire \rf.registers[14][21] ;
 wire \rf.registers[14][22] ;
 wire \rf.registers[14][23] ;
 wire \rf.registers[14][24] ;
 wire \rf.registers[14][25] ;
 wire \rf.registers[14][26] ;
 wire \rf.registers[14][27] ;
 wire \rf.registers[14][28] ;
 wire \rf.registers[14][29] ;
 wire \rf.registers[14][2] ;
 wire \rf.registers[14][30] ;
 wire \rf.registers[14][31] ;
 wire \rf.registers[14][3] ;
 wire \rf.registers[14][4] ;
 wire \rf.registers[14][5] ;
 wire \rf.registers[14][6] ;
 wire \rf.registers[14][7] ;
 wire \rf.registers[14][8] ;
 wire \rf.registers[14][9] ;
 wire \rf.registers[15][0] ;
 wire \rf.registers[15][10] ;
 wire \rf.registers[15][11] ;
 wire \rf.registers[15][12] ;
 wire \rf.registers[15][13] ;
 wire \rf.registers[15][14] ;
 wire \rf.registers[15][15] ;
 wire \rf.registers[15][16] ;
 wire \rf.registers[15][17] ;
 wire \rf.registers[15][18] ;
 wire \rf.registers[15][19] ;
 wire \rf.registers[15][1] ;
 wire \rf.registers[15][20] ;
 wire \rf.registers[15][21] ;
 wire \rf.registers[15][22] ;
 wire \rf.registers[15][23] ;
 wire \rf.registers[15][24] ;
 wire \rf.registers[15][25] ;
 wire \rf.registers[15][26] ;
 wire \rf.registers[15][27] ;
 wire \rf.registers[15][28] ;
 wire \rf.registers[15][29] ;
 wire \rf.registers[15][2] ;
 wire \rf.registers[15][30] ;
 wire \rf.registers[15][31] ;
 wire \rf.registers[15][3] ;
 wire \rf.registers[15][4] ;
 wire \rf.registers[15][5] ;
 wire \rf.registers[15][6] ;
 wire \rf.registers[15][7] ;
 wire \rf.registers[15][8] ;
 wire \rf.registers[15][9] ;
 wire \rf.registers[16][0] ;
 wire \rf.registers[16][10] ;
 wire \rf.registers[16][11] ;
 wire \rf.registers[16][12] ;
 wire \rf.registers[16][13] ;
 wire \rf.registers[16][14] ;
 wire \rf.registers[16][15] ;
 wire \rf.registers[16][16] ;
 wire \rf.registers[16][17] ;
 wire \rf.registers[16][18] ;
 wire \rf.registers[16][19] ;
 wire \rf.registers[16][1] ;
 wire \rf.registers[16][20] ;
 wire \rf.registers[16][21] ;
 wire \rf.registers[16][22] ;
 wire \rf.registers[16][23] ;
 wire \rf.registers[16][24] ;
 wire \rf.registers[16][25] ;
 wire \rf.registers[16][26] ;
 wire \rf.registers[16][27] ;
 wire \rf.registers[16][28] ;
 wire \rf.registers[16][29] ;
 wire \rf.registers[16][2] ;
 wire \rf.registers[16][30] ;
 wire \rf.registers[16][31] ;
 wire \rf.registers[16][3] ;
 wire \rf.registers[16][4] ;
 wire \rf.registers[16][5] ;
 wire \rf.registers[16][6] ;
 wire \rf.registers[16][7] ;
 wire \rf.registers[16][8] ;
 wire \rf.registers[16][9] ;
 wire \rf.registers[17][0] ;
 wire \rf.registers[17][10] ;
 wire \rf.registers[17][11] ;
 wire \rf.registers[17][12] ;
 wire \rf.registers[17][13] ;
 wire \rf.registers[17][14] ;
 wire \rf.registers[17][15] ;
 wire \rf.registers[17][16] ;
 wire \rf.registers[17][17] ;
 wire \rf.registers[17][18] ;
 wire \rf.registers[17][19] ;
 wire \rf.registers[17][1] ;
 wire \rf.registers[17][20] ;
 wire \rf.registers[17][21] ;
 wire \rf.registers[17][22] ;
 wire \rf.registers[17][23] ;
 wire \rf.registers[17][24] ;
 wire \rf.registers[17][25] ;
 wire \rf.registers[17][26] ;
 wire \rf.registers[17][27] ;
 wire \rf.registers[17][28] ;
 wire \rf.registers[17][29] ;
 wire \rf.registers[17][2] ;
 wire \rf.registers[17][30] ;
 wire \rf.registers[17][31] ;
 wire \rf.registers[17][3] ;
 wire \rf.registers[17][4] ;
 wire \rf.registers[17][5] ;
 wire \rf.registers[17][6] ;
 wire \rf.registers[17][7] ;
 wire \rf.registers[17][8] ;
 wire \rf.registers[17][9] ;
 wire \rf.registers[18][0] ;
 wire \rf.registers[18][10] ;
 wire \rf.registers[18][11] ;
 wire \rf.registers[18][12] ;
 wire \rf.registers[18][13] ;
 wire \rf.registers[18][14] ;
 wire \rf.registers[18][15] ;
 wire \rf.registers[18][16] ;
 wire \rf.registers[18][17] ;
 wire \rf.registers[18][18] ;
 wire \rf.registers[18][19] ;
 wire \rf.registers[18][1] ;
 wire \rf.registers[18][20] ;
 wire \rf.registers[18][21] ;
 wire \rf.registers[18][22] ;
 wire \rf.registers[18][23] ;
 wire \rf.registers[18][24] ;
 wire \rf.registers[18][25] ;
 wire \rf.registers[18][26] ;
 wire \rf.registers[18][27] ;
 wire \rf.registers[18][28] ;
 wire \rf.registers[18][29] ;
 wire \rf.registers[18][2] ;
 wire \rf.registers[18][30] ;
 wire \rf.registers[18][31] ;
 wire \rf.registers[18][3] ;
 wire \rf.registers[18][4] ;
 wire \rf.registers[18][5] ;
 wire \rf.registers[18][6] ;
 wire \rf.registers[18][7] ;
 wire \rf.registers[18][8] ;
 wire \rf.registers[18][9] ;
 wire \rf.registers[19][0] ;
 wire \rf.registers[19][10] ;
 wire \rf.registers[19][11] ;
 wire \rf.registers[19][12] ;
 wire \rf.registers[19][13] ;
 wire \rf.registers[19][14] ;
 wire \rf.registers[19][15] ;
 wire \rf.registers[19][16] ;
 wire \rf.registers[19][17] ;
 wire \rf.registers[19][18] ;
 wire \rf.registers[19][19] ;
 wire \rf.registers[19][1] ;
 wire \rf.registers[19][20] ;
 wire \rf.registers[19][21] ;
 wire \rf.registers[19][22] ;
 wire \rf.registers[19][23] ;
 wire \rf.registers[19][24] ;
 wire \rf.registers[19][25] ;
 wire \rf.registers[19][26] ;
 wire \rf.registers[19][27] ;
 wire \rf.registers[19][28] ;
 wire \rf.registers[19][29] ;
 wire \rf.registers[19][2] ;
 wire \rf.registers[19][30] ;
 wire \rf.registers[19][31] ;
 wire \rf.registers[19][3] ;
 wire \rf.registers[19][4] ;
 wire \rf.registers[19][5] ;
 wire \rf.registers[19][6] ;
 wire \rf.registers[19][7] ;
 wire \rf.registers[19][8] ;
 wire \rf.registers[19][9] ;
 wire \rf.registers[1][0] ;
 wire \rf.registers[1][10] ;
 wire \rf.registers[1][11] ;
 wire \rf.registers[1][12] ;
 wire \rf.registers[1][13] ;
 wire \rf.registers[1][14] ;
 wire \rf.registers[1][15] ;
 wire \rf.registers[1][16] ;
 wire \rf.registers[1][17] ;
 wire \rf.registers[1][18] ;
 wire \rf.registers[1][19] ;
 wire \rf.registers[1][1] ;
 wire \rf.registers[1][20] ;
 wire \rf.registers[1][21] ;
 wire \rf.registers[1][22] ;
 wire \rf.registers[1][23] ;
 wire \rf.registers[1][24] ;
 wire \rf.registers[1][25] ;
 wire \rf.registers[1][26] ;
 wire \rf.registers[1][27] ;
 wire \rf.registers[1][28] ;
 wire \rf.registers[1][29] ;
 wire \rf.registers[1][2] ;
 wire \rf.registers[1][30] ;
 wire \rf.registers[1][31] ;
 wire \rf.registers[1][3] ;
 wire \rf.registers[1][4] ;
 wire \rf.registers[1][5] ;
 wire \rf.registers[1][6] ;
 wire \rf.registers[1][7] ;
 wire \rf.registers[1][8] ;
 wire \rf.registers[1][9] ;
 wire \rf.registers[20][0] ;
 wire \rf.registers[20][10] ;
 wire \rf.registers[20][11] ;
 wire \rf.registers[20][12] ;
 wire \rf.registers[20][13] ;
 wire \rf.registers[20][14] ;
 wire \rf.registers[20][15] ;
 wire \rf.registers[20][16] ;
 wire \rf.registers[20][17] ;
 wire \rf.registers[20][18] ;
 wire \rf.registers[20][19] ;
 wire \rf.registers[20][1] ;
 wire \rf.registers[20][20] ;
 wire \rf.registers[20][21] ;
 wire \rf.registers[20][22] ;
 wire \rf.registers[20][23] ;
 wire \rf.registers[20][24] ;
 wire \rf.registers[20][25] ;
 wire \rf.registers[20][26] ;
 wire \rf.registers[20][27] ;
 wire \rf.registers[20][28] ;
 wire \rf.registers[20][29] ;
 wire \rf.registers[20][2] ;
 wire \rf.registers[20][30] ;
 wire \rf.registers[20][31] ;
 wire \rf.registers[20][3] ;
 wire \rf.registers[20][4] ;
 wire \rf.registers[20][5] ;
 wire \rf.registers[20][6] ;
 wire \rf.registers[20][7] ;
 wire \rf.registers[20][8] ;
 wire \rf.registers[20][9] ;
 wire \rf.registers[21][0] ;
 wire \rf.registers[21][10] ;
 wire \rf.registers[21][11] ;
 wire \rf.registers[21][12] ;
 wire \rf.registers[21][13] ;
 wire \rf.registers[21][14] ;
 wire \rf.registers[21][15] ;
 wire \rf.registers[21][16] ;
 wire \rf.registers[21][17] ;
 wire \rf.registers[21][18] ;
 wire \rf.registers[21][19] ;
 wire \rf.registers[21][1] ;
 wire \rf.registers[21][20] ;
 wire \rf.registers[21][21] ;
 wire \rf.registers[21][22] ;
 wire \rf.registers[21][23] ;
 wire \rf.registers[21][24] ;
 wire \rf.registers[21][25] ;
 wire \rf.registers[21][26] ;
 wire \rf.registers[21][27] ;
 wire \rf.registers[21][28] ;
 wire \rf.registers[21][29] ;
 wire \rf.registers[21][2] ;
 wire \rf.registers[21][30] ;
 wire \rf.registers[21][31] ;
 wire \rf.registers[21][3] ;
 wire \rf.registers[21][4] ;
 wire \rf.registers[21][5] ;
 wire \rf.registers[21][6] ;
 wire \rf.registers[21][7] ;
 wire \rf.registers[21][8] ;
 wire \rf.registers[21][9] ;
 wire \rf.registers[22][0] ;
 wire \rf.registers[22][10] ;
 wire \rf.registers[22][11] ;
 wire \rf.registers[22][12] ;
 wire \rf.registers[22][13] ;
 wire \rf.registers[22][14] ;
 wire \rf.registers[22][15] ;
 wire \rf.registers[22][16] ;
 wire \rf.registers[22][17] ;
 wire \rf.registers[22][18] ;
 wire \rf.registers[22][19] ;
 wire \rf.registers[22][1] ;
 wire \rf.registers[22][20] ;
 wire \rf.registers[22][21] ;
 wire \rf.registers[22][22] ;
 wire \rf.registers[22][23] ;
 wire \rf.registers[22][24] ;
 wire \rf.registers[22][25] ;
 wire \rf.registers[22][26] ;
 wire \rf.registers[22][27] ;
 wire \rf.registers[22][28] ;
 wire \rf.registers[22][29] ;
 wire \rf.registers[22][2] ;
 wire \rf.registers[22][30] ;
 wire \rf.registers[22][31] ;
 wire \rf.registers[22][3] ;
 wire \rf.registers[22][4] ;
 wire \rf.registers[22][5] ;
 wire \rf.registers[22][6] ;
 wire \rf.registers[22][7] ;
 wire \rf.registers[22][8] ;
 wire \rf.registers[22][9] ;
 wire \rf.registers[23][0] ;
 wire \rf.registers[23][10] ;
 wire \rf.registers[23][11] ;
 wire \rf.registers[23][12] ;
 wire \rf.registers[23][13] ;
 wire \rf.registers[23][14] ;
 wire \rf.registers[23][15] ;
 wire \rf.registers[23][16] ;
 wire \rf.registers[23][17] ;
 wire \rf.registers[23][18] ;
 wire \rf.registers[23][19] ;
 wire \rf.registers[23][1] ;
 wire \rf.registers[23][20] ;
 wire \rf.registers[23][21] ;
 wire \rf.registers[23][22] ;
 wire \rf.registers[23][23] ;
 wire \rf.registers[23][24] ;
 wire \rf.registers[23][25] ;
 wire \rf.registers[23][26] ;
 wire \rf.registers[23][27] ;
 wire \rf.registers[23][28] ;
 wire \rf.registers[23][29] ;
 wire \rf.registers[23][2] ;
 wire \rf.registers[23][30] ;
 wire \rf.registers[23][31] ;
 wire \rf.registers[23][3] ;
 wire \rf.registers[23][4] ;
 wire \rf.registers[23][5] ;
 wire \rf.registers[23][6] ;
 wire \rf.registers[23][7] ;
 wire \rf.registers[23][8] ;
 wire \rf.registers[23][9] ;
 wire \rf.registers[24][0] ;
 wire \rf.registers[24][10] ;
 wire \rf.registers[24][11] ;
 wire \rf.registers[24][12] ;
 wire \rf.registers[24][13] ;
 wire \rf.registers[24][14] ;
 wire \rf.registers[24][15] ;
 wire \rf.registers[24][16] ;
 wire \rf.registers[24][17] ;
 wire \rf.registers[24][18] ;
 wire \rf.registers[24][19] ;
 wire \rf.registers[24][1] ;
 wire \rf.registers[24][20] ;
 wire \rf.registers[24][21] ;
 wire \rf.registers[24][22] ;
 wire \rf.registers[24][23] ;
 wire \rf.registers[24][24] ;
 wire \rf.registers[24][25] ;
 wire \rf.registers[24][26] ;
 wire \rf.registers[24][27] ;
 wire \rf.registers[24][28] ;
 wire \rf.registers[24][29] ;
 wire \rf.registers[24][2] ;
 wire \rf.registers[24][30] ;
 wire \rf.registers[24][31] ;
 wire \rf.registers[24][3] ;
 wire \rf.registers[24][4] ;
 wire \rf.registers[24][5] ;
 wire \rf.registers[24][6] ;
 wire \rf.registers[24][7] ;
 wire \rf.registers[24][8] ;
 wire \rf.registers[24][9] ;
 wire \rf.registers[25][0] ;
 wire \rf.registers[25][10] ;
 wire \rf.registers[25][11] ;
 wire \rf.registers[25][12] ;
 wire \rf.registers[25][13] ;
 wire \rf.registers[25][14] ;
 wire \rf.registers[25][15] ;
 wire \rf.registers[25][16] ;
 wire \rf.registers[25][17] ;
 wire \rf.registers[25][18] ;
 wire \rf.registers[25][19] ;
 wire \rf.registers[25][1] ;
 wire \rf.registers[25][20] ;
 wire \rf.registers[25][21] ;
 wire \rf.registers[25][22] ;
 wire \rf.registers[25][23] ;
 wire \rf.registers[25][24] ;
 wire \rf.registers[25][25] ;
 wire \rf.registers[25][26] ;
 wire \rf.registers[25][27] ;
 wire \rf.registers[25][28] ;
 wire \rf.registers[25][29] ;
 wire \rf.registers[25][2] ;
 wire \rf.registers[25][30] ;
 wire \rf.registers[25][31] ;
 wire \rf.registers[25][3] ;
 wire \rf.registers[25][4] ;
 wire \rf.registers[25][5] ;
 wire \rf.registers[25][6] ;
 wire \rf.registers[25][7] ;
 wire \rf.registers[25][8] ;
 wire \rf.registers[25][9] ;
 wire \rf.registers[26][0] ;
 wire \rf.registers[26][10] ;
 wire \rf.registers[26][11] ;
 wire \rf.registers[26][12] ;
 wire \rf.registers[26][13] ;
 wire \rf.registers[26][14] ;
 wire \rf.registers[26][15] ;
 wire \rf.registers[26][16] ;
 wire \rf.registers[26][17] ;
 wire \rf.registers[26][18] ;
 wire \rf.registers[26][19] ;
 wire \rf.registers[26][1] ;
 wire \rf.registers[26][20] ;
 wire \rf.registers[26][21] ;
 wire \rf.registers[26][22] ;
 wire \rf.registers[26][23] ;
 wire \rf.registers[26][24] ;
 wire \rf.registers[26][25] ;
 wire \rf.registers[26][26] ;
 wire \rf.registers[26][27] ;
 wire \rf.registers[26][28] ;
 wire \rf.registers[26][29] ;
 wire \rf.registers[26][2] ;
 wire \rf.registers[26][30] ;
 wire \rf.registers[26][31] ;
 wire \rf.registers[26][3] ;
 wire \rf.registers[26][4] ;
 wire \rf.registers[26][5] ;
 wire \rf.registers[26][6] ;
 wire \rf.registers[26][7] ;
 wire \rf.registers[26][8] ;
 wire \rf.registers[26][9] ;
 wire \rf.registers[27][0] ;
 wire \rf.registers[27][10] ;
 wire \rf.registers[27][11] ;
 wire \rf.registers[27][12] ;
 wire \rf.registers[27][13] ;
 wire \rf.registers[27][14] ;
 wire \rf.registers[27][15] ;
 wire \rf.registers[27][16] ;
 wire \rf.registers[27][17] ;
 wire \rf.registers[27][18] ;
 wire \rf.registers[27][19] ;
 wire \rf.registers[27][1] ;
 wire \rf.registers[27][20] ;
 wire \rf.registers[27][21] ;
 wire \rf.registers[27][22] ;
 wire \rf.registers[27][23] ;
 wire \rf.registers[27][24] ;
 wire \rf.registers[27][25] ;
 wire \rf.registers[27][26] ;
 wire \rf.registers[27][27] ;
 wire \rf.registers[27][28] ;
 wire \rf.registers[27][29] ;
 wire \rf.registers[27][2] ;
 wire \rf.registers[27][30] ;
 wire \rf.registers[27][31] ;
 wire \rf.registers[27][3] ;
 wire \rf.registers[27][4] ;
 wire \rf.registers[27][5] ;
 wire \rf.registers[27][6] ;
 wire \rf.registers[27][7] ;
 wire \rf.registers[27][8] ;
 wire \rf.registers[27][9] ;
 wire \rf.registers[28][0] ;
 wire \rf.registers[28][10] ;
 wire \rf.registers[28][11] ;
 wire \rf.registers[28][12] ;
 wire \rf.registers[28][13] ;
 wire \rf.registers[28][14] ;
 wire \rf.registers[28][15] ;
 wire \rf.registers[28][16] ;
 wire \rf.registers[28][17] ;
 wire \rf.registers[28][18] ;
 wire \rf.registers[28][19] ;
 wire \rf.registers[28][1] ;
 wire \rf.registers[28][20] ;
 wire \rf.registers[28][21] ;
 wire \rf.registers[28][22] ;
 wire \rf.registers[28][23] ;
 wire \rf.registers[28][24] ;
 wire \rf.registers[28][25] ;
 wire \rf.registers[28][26] ;
 wire \rf.registers[28][27] ;
 wire \rf.registers[28][28] ;
 wire \rf.registers[28][29] ;
 wire \rf.registers[28][2] ;
 wire \rf.registers[28][30] ;
 wire \rf.registers[28][31] ;
 wire \rf.registers[28][3] ;
 wire \rf.registers[28][4] ;
 wire \rf.registers[28][5] ;
 wire \rf.registers[28][6] ;
 wire \rf.registers[28][7] ;
 wire \rf.registers[28][8] ;
 wire \rf.registers[28][9] ;
 wire \rf.registers[29][0] ;
 wire \rf.registers[29][10] ;
 wire \rf.registers[29][11] ;
 wire \rf.registers[29][12] ;
 wire \rf.registers[29][13] ;
 wire \rf.registers[29][14] ;
 wire \rf.registers[29][15] ;
 wire \rf.registers[29][16] ;
 wire \rf.registers[29][17] ;
 wire \rf.registers[29][18] ;
 wire \rf.registers[29][19] ;
 wire \rf.registers[29][1] ;
 wire \rf.registers[29][20] ;
 wire \rf.registers[29][21] ;
 wire \rf.registers[29][22] ;
 wire \rf.registers[29][23] ;
 wire \rf.registers[29][24] ;
 wire \rf.registers[29][25] ;
 wire \rf.registers[29][26] ;
 wire \rf.registers[29][27] ;
 wire \rf.registers[29][28] ;
 wire \rf.registers[29][29] ;
 wire \rf.registers[29][2] ;
 wire \rf.registers[29][30] ;
 wire \rf.registers[29][31] ;
 wire \rf.registers[29][3] ;
 wire \rf.registers[29][4] ;
 wire \rf.registers[29][5] ;
 wire \rf.registers[29][6] ;
 wire \rf.registers[29][7] ;
 wire \rf.registers[29][8] ;
 wire \rf.registers[29][9] ;
 wire \rf.registers[2][0] ;
 wire \rf.registers[2][10] ;
 wire \rf.registers[2][11] ;
 wire \rf.registers[2][12] ;
 wire \rf.registers[2][13] ;
 wire \rf.registers[2][14] ;
 wire \rf.registers[2][15] ;
 wire \rf.registers[2][16] ;
 wire \rf.registers[2][17] ;
 wire \rf.registers[2][18] ;
 wire \rf.registers[2][19] ;
 wire \rf.registers[2][1] ;
 wire \rf.registers[2][20] ;
 wire \rf.registers[2][21] ;
 wire \rf.registers[2][22] ;
 wire \rf.registers[2][23] ;
 wire \rf.registers[2][24] ;
 wire \rf.registers[2][25] ;
 wire \rf.registers[2][26] ;
 wire \rf.registers[2][27] ;
 wire \rf.registers[2][28] ;
 wire \rf.registers[2][29] ;
 wire \rf.registers[2][2] ;
 wire \rf.registers[2][30] ;
 wire \rf.registers[2][31] ;
 wire \rf.registers[2][3] ;
 wire \rf.registers[2][4] ;
 wire \rf.registers[2][5] ;
 wire \rf.registers[2][6] ;
 wire \rf.registers[2][7] ;
 wire \rf.registers[2][8] ;
 wire \rf.registers[2][9] ;
 wire \rf.registers[30][0] ;
 wire \rf.registers[30][10] ;
 wire \rf.registers[30][11] ;
 wire \rf.registers[30][12] ;
 wire \rf.registers[30][13] ;
 wire \rf.registers[30][14] ;
 wire \rf.registers[30][15] ;
 wire \rf.registers[30][16] ;
 wire \rf.registers[30][17] ;
 wire \rf.registers[30][18] ;
 wire \rf.registers[30][19] ;
 wire \rf.registers[30][1] ;
 wire \rf.registers[30][20] ;
 wire \rf.registers[30][21] ;
 wire \rf.registers[30][22] ;
 wire \rf.registers[30][23] ;
 wire \rf.registers[30][24] ;
 wire \rf.registers[30][25] ;
 wire \rf.registers[30][26] ;
 wire \rf.registers[30][27] ;
 wire \rf.registers[30][28] ;
 wire \rf.registers[30][29] ;
 wire \rf.registers[30][2] ;
 wire \rf.registers[30][30] ;
 wire \rf.registers[30][31] ;
 wire \rf.registers[30][3] ;
 wire \rf.registers[30][4] ;
 wire \rf.registers[30][5] ;
 wire \rf.registers[30][6] ;
 wire \rf.registers[30][7] ;
 wire \rf.registers[30][8] ;
 wire \rf.registers[30][9] ;
 wire \rf.registers[31][0] ;
 wire \rf.registers[31][10] ;
 wire \rf.registers[31][11] ;
 wire \rf.registers[31][12] ;
 wire \rf.registers[31][13] ;
 wire \rf.registers[31][14] ;
 wire \rf.registers[31][15] ;
 wire \rf.registers[31][16] ;
 wire \rf.registers[31][17] ;
 wire \rf.registers[31][18] ;
 wire \rf.registers[31][19] ;
 wire \rf.registers[31][1] ;
 wire \rf.registers[31][20] ;
 wire \rf.registers[31][21] ;
 wire \rf.registers[31][22] ;
 wire \rf.registers[31][23] ;
 wire \rf.registers[31][24] ;
 wire \rf.registers[31][25] ;
 wire \rf.registers[31][26] ;
 wire \rf.registers[31][27] ;
 wire \rf.registers[31][28] ;
 wire \rf.registers[31][29] ;
 wire \rf.registers[31][2] ;
 wire \rf.registers[31][30] ;
 wire \rf.registers[31][31] ;
 wire \rf.registers[31][3] ;
 wire \rf.registers[31][4] ;
 wire \rf.registers[31][5] ;
 wire \rf.registers[31][6] ;
 wire \rf.registers[31][7] ;
 wire \rf.registers[31][8] ;
 wire \rf.registers[31][9] ;
 wire \rf.registers[3][0] ;
 wire \rf.registers[3][10] ;
 wire \rf.registers[3][11] ;
 wire \rf.registers[3][12] ;
 wire \rf.registers[3][13] ;
 wire \rf.registers[3][14] ;
 wire \rf.registers[3][15] ;
 wire \rf.registers[3][16] ;
 wire \rf.registers[3][17] ;
 wire \rf.registers[3][18] ;
 wire \rf.registers[3][19] ;
 wire \rf.registers[3][1] ;
 wire \rf.registers[3][20] ;
 wire \rf.registers[3][21] ;
 wire \rf.registers[3][22] ;
 wire \rf.registers[3][23] ;
 wire \rf.registers[3][24] ;
 wire \rf.registers[3][25] ;
 wire \rf.registers[3][26] ;
 wire \rf.registers[3][27] ;
 wire \rf.registers[3][28] ;
 wire \rf.registers[3][29] ;
 wire \rf.registers[3][2] ;
 wire \rf.registers[3][30] ;
 wire \rf.registers[3][31] ;
 wire \rf.registers[3][3] ;
 wire \rf.registers[3][4] ;
 wire \rf.registers[3][5] ;
 wire \rf.registers[3][6] ;
 wire \rf.registers[3][7] ;
 wire \rf.registers[3][8] ;
 wire \rf.registers[3][9] ;
 wire \rf.registers[4][0] ;
 wire \rf.registers[4][10] ;
 wire \rf.registers[4][11] ;
 wire \rf.registers[4][12] ;
 wire \rf.registers[4][13] ;
 wire \rf.registers[4][14] ;
 wire \rf.registers[4][15] ;
 wire \rf.registers[4][16] ;
 wire \rf.registers[4][17] ;
 wire \rf.registers[4][18] ;
 wire \rf.registers[4][19] ;
 wire \rf.registers[4][1] ;
 wire \rf.registers[4][20] ;
 wire \rf.registers[4][21] ;
 wire \rf.registers[4][22] ;
 wire \rf.registers[4][23] ;
 wire \rf.registers[4][24] ;
 wire \rf.registers[4][25] ;
 wire \rf.registers[4][26] ;
 wire \rf.registers[4][27] ;
 wire \rf.registers[4][28] ;
 wire \rf.registers[4][29] ;
 wire \rf.registers[4][2] ;
 wire \rf.registers[4][30] ;
 wire \rf.registers[4][31] ;
 wire \rf.registers[4][3] ;
 wire \rf.registers[4][4] ;
 wire \rf.registers[4][5] ;
 wire \rf.registers[4][6] ;
 wire \rf.registers[4][7] ;
 wire \rf.registers[4][8] ;
 wire \rf.registers[4][9] ;
 wire \rf.registers[5][0] ;
 wire \rf.registers[5][10] ;
 wire \rf.registers[5][11] ;
 wire \rf.registers[5][12] ;
 wire \rf.registers[5][13] ;
 wire \rf.registers[5][14] ;
 wire \rf.registers[5][15] ;
 wire \rf.registers[5][16] ;
 wire \rf.registers[5][17] ;
 wire \rf.registers[5][18] ;
 wire \rf.registers[5][19] ;
 wire \rf.registers[5][1] ;
 wire \rf.registers[5][20] ;
 wire \rf.registers[5][21] ;
 wire \rf.registers[5][22] ;
 wire \rf.registers[5][23] ;
 wire \rf.registers[5][24] ;
 wire \rf.registers[5][25] ;
 wire \rf.registers[5][26] ;
 wire \rf.registers[5][27] ;
 wire \rf.registers[5][28] ;
 wire \rf.registers[5][29] ;
 wire \rf.registers[5][2] ;
 wire \rf.registers[5][30] ;
 wire \rf.registers[5][31] ;
 wire \rf.registers[5][3] ;
 wire \rf.registers[5][4] ;
 wire \rf.registers[5][5] ;
 wire \rf.registers[5][6] ;
 wire \rf.registers[5][7] ;
 wire \rf.registers[5][8] ;
 wire \rf.registers[5][9] ;
 wire \rf.registers[6][0] ;
 wire \rf.registers[6][10] ;
 wire \rf.registers[6][11] ;
 wire \rf.registers[6][12] ;
 wire \rf.registers[6][13] ;
 wire \rf.registers[6][14] ;
 wire \rf.registers[6][15] ;
 wire \rf.registers[6][16] ;
 wire \rf.registers[6][17] ;
 wire \rf.registers[6][18] ;
 wire \rf.registers[6][19] ;
 wire \rf.registers[6][1] ;
 wire \rf.registers[6][20] ;
 wire \rf.registers[6][21] ;
 wire \rf.registers[6][22] ;
 wire \rf.registers[6][23] ;
 wire \rf.registers[6][24] ;
 wire \rf.registers[6][25] ;
 wire \rf.registers[6][26] ;
 wire \rf.registers[6][27] ;
 wire \rf.registers[6][28] ;
 wire \rf.registers[6][29] ;
 wire \rf.registers[6][2] ;
 wire \rf.registers[6][30] ;
 wire \rf.registers[6][31] ;
 wire \rf.registers[6][3] ;
 wire \rf.registers[6][4] ;
 wire \rf.registers[6][5] ;
 wire \rf.registers[6][6] ;
 wire \rf.registers[6][7] ;
 wire \rf.registers[6][8] ;
 wire \rf.registers[6][9] ;
 wire \rf.registers[7][0] ;
 wire \rf.registers[7][10] ;
 wire \rf.registers[7][11] ;
 wire \rf.registers[7][12] ;
 wire \rf.registers[7][13] ;
 wire \rf.registers[7][14] ;
 wire \rf.registers[7][15] ;
 wire \rf.registers[7][16] ;
 wire \rf.registers[7][17] ;
 wire \rf.registers[7][18] ;
 wire \rf.registers[7][19] ;
 wire \rf.registers[7][1] ;
 wire \rf.registers[7][20] ;
 wire \rf.registers[7][21] ;
 wire \rf.registers[7][22] ;
 wire \rf.registers[7][23] ;
 wire \rf.registers[7][24] ;
 wire \rf.registers[7][25] ;
 wire \rf.registers[7][26] ;
 wire \rf.registers[7][27] ;
 wire \rf.registers[7][28] ;
 wire \rf.registers[7][29] ;
 wire \rf.registers[7][2] ;
 wire \rf.registers[7][30] ;
 wire \rf.registers[7][31] ;
 wire \rf.registers[7][3] ;
 wire \rf.registers[7][4] ;
 wire \rf.registers[7][5] ;
 wire \rf.registers[7][6] ;
 wire \rf.registers[7][7] ;
 wire \rf.registers[7][8] ;
 wire \rf.registers[7][9] ;
 wire \rf.registers[8][0] ;
 wire \rf.registers[8][10] ;
 wire \rf.registers[8][11] ;
 wire \rf.registers[8][12] ;
 wire \rf.registers[8][13] ;
 wire \rf.registers[8][14] ;
 wire \rf.registers[8][15] ;
 wire \rf.registers[8][16] ;
 wire \rf.registers[8][17] ;
 wire \rf.registers[8][18] ;
 wire \rf.registers[8][19] ;
 wire \rf.registers[8][1] ;
 wire \rf.registers[8][20] ;
 wire \rf.registers[8][21] ;
 wire \rf.registers[8][22] ;
 wire \rf.registers[8][23] ;
 wire \rf.registers[8][24] ;
 wire \rf.registers[8][25] ;
 wire \rf.registers[8][26] ;
 wire \rf.registers[8][27] ;
 wire \rf.registers[8][28] ;
 wire \rf.registers[8][29] ;
 wire \rf.registers[8][2] ;
 wire \rf.registers[8][30] ;
 wire \rf.registers[8][31] ;
 wire \rf.registers[8][3] ;
 wire \rf.registers[8][4] ;
 wire \rf.registers[8][5] ;
 wire \rf.registers[8][6] ;
 wire \rf.registers[8][7] ;
 wire \rf.registers[8][8] ;
 wire \rf.registers[8][9] ;
 wire \rf.registers[9][0] ;
 wire \rf.registers[9][10] ;
 wire \rf.registers[9][11] ;
 wire \rf.registers[9][12] ;
 wire \rf.registers[9][13] ;
 wire \rf.registers[9][14] ;
 wire \rf.registers[9][15] ;
 wire \rf.registers[9][16] ;
 wire \rf.registers[9][17] ;
 wire \rf.registers[9][18] ;
 wire \rf.registers[9][19] ;
 wire \rf.registers[9][1] ;
 wire \rf.registers[9][20] ;
 wire \rf.registers[9][21] ;
 wire \rf.registers[9][22] ;
 wire \rf.registers[9][23] ;
 wire \rf.registers[9][24] ;
 wire \rf.registers[9][25] ;
 wire \rf.registers[9][26] ;
 wire \rf.registers[9][27] ;
 wire \rf.registers[9][28] ;
 wire \rf.registers[9][29] ;
 wire \rf.registers[9][2] ;
 wire \rf.registers[9][30] ;
 wire \rf.registers[9][31] ;
 wire \rf.registers[9][3] ;
 wire \rf.registers[9][4] ;
 wire \rf.registers[9][5] ;
 wire \rf.registers[9][6] ;
 wire \rf.registers[9][7] ;
 wire \rf.registers[9][8] ;
 wire \rf.registers[9][9] ;

 sky130_fd_sc_hd__inv_2 _4268_ (.A(A2[4]),
    .Y(_1024_));
 sky130_fd_sc_hd__buf_1 _4269_ (.A(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__buf_1 _4270_ (.A(A2[0]),
    .X(_1026_));
 sky130_fd_sc_hd__buf_1 _4271_ (.A(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__buf_1 _4272_ (.A(A2[1]),
    .X(_1028_));
 sky130_fd_sc_hd__buf_1 _4273_ (.A(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__mux4_2 _4274_ (.A0(\rf.registers[20][4] ),
    .A1(\rf.registers[21][4] ),
    .A2(\rf.registers[22][4] ),
    .A3(\rf.registers[23][4] ),
    .S0(_1027_),
    .S1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__mux4_2 _4275_ (.A0(\rf.registers[16][4] ),
    .A1(\rf.registers[17][4] ),
    .A2(\rf.registers[18][4] ),
    .A3(\rf.registers[19][4] ),
    .S0(_1027_),
    .S1(_1029_),
    .X(_1031_));
 sky130_fd_sc_hd__mux4_2 _4276_ (.A0(\rf.registers[28][4] ),
    .A1(\rf.registers[29][4] ),
    .A2(\rf.registers[30][4] ),
    .A3(\rf.registers[31][4] ),
    .S0(_1027_),
    .S1(_1029_),
    .X(_1032_));
 sky130_fd_sc_hd__mux4_2 _4277_ (.A0(\rf.registers[24][4] ),
    .A1(\rf.registers[25][4] ),
    .A2(\rf.registers[26][4] ),
    .A3(\rf.registers[27][4] ),
    .S0(_1027_),
    .S1(_1029_),
    .X(_1033_));
 sky130_fd_sc_hd__inv_2 _4278_ (.A(A2[2]),
    .Y(_1034_));
 sky130_fd_sc_hd__buf_1 _4279_ (.A(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__buf_1 _4280_ (.A(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__buf_1 _4281_ (.A(A2[3]),
    .X(_1037_));
 sky130_fd_sc_hd__buf_1 _4282_ (.A(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__mux4_2 _4283_ (.A0(_1030_),
    .A1(_1031_),
    .A2(_1032_),
    .A3(_1033_),
    .S0(_1036_),
    .S1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__buf_1 _4284_ (.A(_1034_),
    .X(_1040_));
 sky130_fd_sc_hd__buf_1 _4285_ (.A(A2[0]),
    .X(_1041_));
 sky130_fd_sc_hd__buf_1 _4286_ (.A(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__buf_1 _4287_ (.A(A2[1]),
    .X(_1043_));
 sky130_fd_sc_hd__buf_1 _4288_ (.A(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__mux4_2 _4289_ (.A0(\rf.registers[4][4] ),
    .A1(\rf.registers[5][4] ),
    .A2(\rf.registers[6][4] ),
    .A3(\rf.registers[7][4] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__or2_2 _4290_ (.A(_1040_),
    .B(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__buf_1 _4291_ (.A(A2[2]),
    .X(_1047_));
 sky130_fd_sc_hd__buf_1 _4292_ (.A(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__mux4_2 _4293_ (.A0(\rf.registers[0][4] ),
    .A1(\rf.registers[1][4] ),
    .A2(\rf.registers[2][4] ),
    .A3(\rf.registers[3][4] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1049_));
 sky130_fd_sc_hd__inv_2 _4294_ (.A(A2[3]),
    .Y(_1050_));
 sky130_fd_sc_hd__o21a_2 _4295_ (.A1(_1048_),
    .A2(_1049_),
    .B1(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__buf_1 _4296_ (.A(_1041_),
    .X(_1052_));
 sky130_fd_sc_hd__buf_1 _4297_ (.A(_1043_),
    .X(_1053_));
 sky130_fd_sc_hd__mux4_2 _4298_ (.A0(\rf.registers[8][4] ),
    .A1(\rf.registers[9][4] ),
    .A2(\rf.registers[10][4] ),
    .A3(\rf.registers[11][4] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__mux4_2 _4299_ (.A0(\rf.registers[12][4] ),
    .A1(\rf.registers[13][4] ),
    .A2(\rf.registers[14][4] ),
    .A3(\rf.registers[15][4] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1055_));
 sky130_fd_sc_hd__mux2_2 _4300_ (.A0(_1054_),
    .A1(_1055_),
    .S(_1047_),
    .X(_1056_));
 sky130_fd_sc_hd__buf_1 _4301_ (.A(A2[4]),
    .X(_1057_));
 sky130_fd_sc_hd__a221o_2 _4302_ (.A1(_1046_),
    .A2(_1051_),
    .B1(_1056_),
    .B2(_1038_),
    .C1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__o21ai_2 _4303_ (.A1(_1025_),
    .A2(_1039_),
    .B1(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__buf_1 _4304_ (.A(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__buf_1 _4305_ (.A(A2[1]),
    .X(_1061_));
 sky130_fd_sc_hd__mux4_2 _4306_ (.A0(\rf.registers[20][5] ),
    .A1(\rf.registers[21][5] ),
    .A2(\rf.registers[22][5] ),
    .A3(\rf.registers[23][5] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__mux4_2 _4307_ (.A0(\rf.registers[16][5] ),
    .A1(\rf.registers[17][5] ),
    .A2(\rf.registers[18][5] ),
    .A3(\rf.registers[19][5] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_2 _4308_ (.A0(_1062_),
    .A1(_1063_),
    .S(_1035_),
    .X(_1064_));
 sky130_fd_sc_hd__buf_1 _4309_ (.A(A2[0]),
    .X(_1065_));
 sky130_fd_sc_hd__buf_1 _4310_ (.A(A2[1]),
    .X(_1066_));
 sky130_fd_sc_hd__mux4_2 _4311_ (.A0(\rf.registers[28][5] ),
    .A1(\rf.registers[29][5] ),
    .A2(\rf.registers[30][5] ),
    .A3(\rf.registers[31][5] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__mux4_2 _4312_ (.A0(\rf.registers[24][5] ),
    .A1(\rf.registers[25][5] ),
    .A2(\rf.registers[26][5] ),
    .A3(\rf.registers[27][5] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_2 _4313_ (.A0(_1067_),
    .A1(_1068_),
    .S(_1035_),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_2 _4314_ (.A0(_1064_),
    .A1(_1069_),
    .S(_1037_),
    .X(_1070_));
 sky130_fd_sc_hd__buf_1 _4315_ (.A(_1037_),
    .X(_1071_));
 sky130_fd_sc_hd__buf_1 _4316_ (.A(_1041_),
    .X(_1072_));
 sky130_fd_sc_hd__buf_1 _4317_ (.A(_1043_),
    .X(_1073_));
 sky130_fd_sc_hd__mux4_2 _4318_ (.A0(\rf.registers[8][5] ),
    .A1(\rf.registers[9][5] ),
    .A2(\rf.registers[10][5] ),
    .A3(\rf.registers[11][5] ),
    .S0(_1072_),
    .S1(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__mux4_2 _4319_ (.A0(\rf.registers[12][5] ),
    .A1(\rf.registers[13][5] ),
    .A2(\rf.registers[14][5] ),
    .A3(\rf.registers[15][5] ),
    .S0(_1072_),
    .S1(_1073_),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_2 _4320_ (.A0(_1074_),
    .A1(_1075_),
    .S(_1048_),
    .X(_1076_));
 sky130_fd_sc_hd__nand2_2 _4321_ (.A(_1071_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__buf_1 _4322_ (.A(_1050_),
    .X(_1078_));
 sky130_fd_sc_hd__mux4_2 _4323_ (.A0(\rf.registers[4][5] ),
    .A1(\rf.registers[5][5] ),
    .A2(\rf.registers[6][5] ),
    .A3(\rf.registers[7][5] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1079_));
 sky130_fd_sc_hd__mux4_2 _4324_ (.A0(\rf.registers[0][5] ),
    .A1(\rf.registers[1][5] ),
    .A2(\rf.registers[2][5] ),
    .A3(\rf.registers[3][5] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1080_));
 sky130_fd_sc_hd__mux2_2 _4325_ (.A0(_1079_),
    .A1(_1080_),
    .S(_1040_),
    .X(_1081_));
 sky130_fd_sc_hd__a21oi_2 _4326_ (.A1(_1078_),
    .A2(_1081_),
    .B1(_1057_),
    .Y(_1082_));
 sky130_fd_sc_hd__a2bb2o_2 _4327_ (.A1_N(_1025_),
    .A2_N(_1070_),
    .B1(_1077_),
    .B2(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__nand2_2 _4328_ (.A(opcode[1]),
    .B(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__nor2_2 _4329_ (.A(opcode[0]),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__and2_2 _4330_ (.A(_1060_),
    .B(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__buf_1 _4331_ (.A(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__buf_1 _4332_ (.A(_1050_),
    .X(_1088_));
 sky130_fd_sc_hd__buf_1 _4333_ (.A(_1041_),
    .X(_1089_));
 sky130_fd_sc_hd__buf_1 _4334_ (.A(_1043_),
    .X(_1090_));
 sky130_fd_sc_hd__mux4_2 _4335_ (.A0(\rf.registers[20][3] ),
    .A1(\rf.registers[21][3] ),
    .A2(\rf.registers[22][3] ),
    .A3(\rf.registers[23][3] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__mux4_2 _4336_ (.A0(\rf.registers[16][3] ),
    .A1(\rf.registers[17][3] ),
    .A2(\rf.registers[18][3] ),
    .A3(\rf.registers[19][3] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_2 _4337_ (.A0(_1091_),
    .A1(_1092_),
    .S(_1040_),
    .X(_1093_));
 sky130_fd_sc_hd__nand2_2 _4338_ (.A(_1088_),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__mux4_2 _4339_ (.A0(\rf.registers[28][3] ),
    .A1(\rf.registers[29][3] ),
    .A2(\rf.registers[30][3] ),
    .A3(\rf.registers[31][3] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1095_));
 sky130_fd_sc_hd__mux4_2 _4340_ (.A0(\rf.registers[24][3] ),
    .A1(\rf.registers[25][3] ),
    .A2(\rf.registers[26][3] ),
    .A3(\rf.registers[27][3] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_2 _4341_ (.A0(_1095_),
    .A1(_1096_),
    .S(_1040_),
    .X(_1097_));
 sky130_fd_sc_hd__nand2_2 _4342_ (.A(_1038_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__mux4_2 _4343_ (.A0(\rf.registers[8][3] ),
    .A1(\rf.registers[9][3] ),
    .A2(\rf.registers[10][3] ),
    .A3(\rf.registers[11][3] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1099_));
 sky130_fd_sc_hd__mux4_2 _4344_ (.A0(\rf.registers[12][3] ),
    .A1(\rf.registers[13][3] ),
    .A2(\rf.registers[14][3] ),
    .A3(\rf.registers[15][3] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_2 _4345_ (.A0(_1099_),
    .A1(_1100_),
    .S(_1048_),
    .X(_1101_));
 sky130_fd_sc_hd__nand2_2 _4346_ (.A(_1071_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__mux4_2 _4347_ (.A0(\rf.registers[4][3] ),
    .A1(\rf.registers[5][3] ),
    .A2(\rf.registers[6][3] ),
    .A3(\rf.registers[7][3] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1103_));
 sky130_fd_sc_hd__buf_1 _4348_ (.A(_1041_),
    .X(_1104_));
 sky130_fd_sc_hd__buf_1 _4349_ (.A(_1043_),
    .X(_1105_));
 sky130_fd_sc_hd__mux4_2 _4350_ (.A0(\rf.registers[0][3] ),
    .A1(\rf.registers[1][3] ),
    .A2(\rf.registers[2][3] ),
    .A3(\rf.registers[3][3] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__buf_1 _4351_ (.A(_1034_),
    .X(_1107_));
 sky130_fd_sc_hd__mux2_2 _4352_ (.A0(_1103_),
    .A1(_1106_),
    .S(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__a21oi_2 _4353_ (.A1(_1088_),
    .A2(_1108_),
    .B1(A2[4]),
    .Y(_1109_));
 sky130_fd_sc_hd__a32o_2 _4354_ (.A1(_1057_),
    .A2(_1094_),
    .A3(_1098_),
    .B1(_1102_),
    .B2(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__buf_1 _4355_ (.A(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__mux4_2 _4356_ (.A0(\rf.registers[24][2] ),
    .A1(\rf.registers[25][2] ),
    .A2(\rf.registers[26][2] ),
    .A3(\rf.registers[27][2] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1112_));
 sky130_fd_sc_hd__mux4_2 _4357_ (.A0(\rf.registers[28][2] ),
    .A1(\rf.registers[29][2] ),
    .A2(\rf.registers[30][2] ),
    .A3(\rf.registers[31][2] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1113_));
 sky130_fd_sc_hd__mux4_2 _4358_ (.A0(\rf.registers[16][2] ),
    .A1(\rf.registers[17][2] ),
    .A2(\rf.registers[18][2] ),
    .A3(\rf.registers[19][2] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1114_));
 sky130_fd_sc_hd__mux4_2 _4359_ (.A0(\rf.registers[20][2] ),
    .A1(\rf.registers[21][2] ),
    .A2(\rf.registers[22][2] ),
    .A3(\rf.registers[23][2] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1115_));
 sky130_fd_sc_hd__mux4_2 _4360_ (.A0(_1112_),
    .A1(_1113_),
    .A2(_1114_),
    .A3(_1115_),
    .S0(_1047_),
    .S1(_1050_),
    .X(_1116_));
 sky130_fd_sc_hd__mux4_2 _4361_ (.A0(\rf.registers[4][2] ),
    .A1(\rf.registers[5][2] ),
    .A2(\rf.registers[6][2] ),
    .A3(\rf.registers[7][2] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1117_));
 sky130_fd_sc_hd__or2_2 _4362_ (.A(_1107_),
    .B(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__mux4_2 _4363_ (.A0(\rf.registers[0][2] ),
    .A1(\rf.registers[1][2] ),
    .A2(\rf.registers[2][2] ),
    .A3(\rf.registers[3][2] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1119_));
 sky130_fd_sc_hd__o21a_2 _4364_ (.A1(_1047_),
    .A2(_1119_),
    .B1(_1050_),
    .X(_1120_));
 sky130_fd_sc_hd__mux4_2 _4365_ (.A0(\rf.registers[8][2] ),
    .A1(\rf.registers[9][2] ),
    .A2(\rf.registers[10][2] ),
    .A3(\rf.registers[11][2] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1121_));
 sky130_fd_sc_hd__mux4_2 _4366_ (.A0(\rf.registers[12][2] ),
    .A1(\rf.registers[13][2] ),
    .A2(\rf.registers[14][2] ),
    .A3(\rf.registers[15][2] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1122_));
 sky130_fd_sc_hd__mux2_2 _4367_ (.A0(_1121_),
    .A1(_1122_),
    .S(_1047_),
    .X(_1123_));
 sky130_fd_sc_hd__a221o_2 _4368_ (.A1(_1118_),
    .A2(_1120_),
    .B1(_1123_),
    .B2(_1037_),
    .C1(A2[4]),
    .X(_1124_));
 sky130_fd_sc_hd__o21ai_2 _4369_ (.A1(_1024_),
    .A2(_1116_),
    .B1(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__buf_1 _4370_ (.A(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__and2_2 _4371_ (.A(_1111_),
    .B(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__nand2_2 _4372_ (.A(_1087_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__mux4_2 _4373_ (.A0(\rf.registers[20][1] ),
    .A1(\rf.registers[21][1] ),
    .A2(\rf.registers[22][1] ),
    .A3(\rf.registers[23][1] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1129_));
 sky130_fd_sc_hd__mux4_2 _4374_ (.A0(\rf.registers[16][1] ),
    .A1(\rf.registers[17][1] ),
    .A2(\rf.registers[18][1] ),
    .A3(\rf.registers[19][1] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_2 _4375_ (.A0(_1129_),
    .A1(_1130_),
    .S(_1035_),
    .X(_1131_));
 sky130_fd_sc_hd__mux4_2 _4376_ (.A0(\rf.registers[28][1] ),
    .A1(\rf.registers[29][1] ),
    .A2(\rf.registers[30][1] ),
    .A3(\rf.registers[31][1] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1132_));
 sky130_fd_sc_hd__mux4_2 _4377_ (.A0(\rf.registers[24][1] ),
    .A1(\rf.registers[25][1] ),
    .A2(\rf.registers[26][1] ),
    .A3(\rf.registers[27][1] ),
    .S0(_1041_),
    .S1(_1043_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_2 _4378_ (.A0(_1132_),
    .A1(_1133_),
    .S(_1035_),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_2 _4379_ (.A0(_1131_),
    .A1(_1134_),
    .S(_1037_),
    .X(_1135_));
 sky130_fd_sc_hd__mux4_2 _4380_ (.A0(\rf.registers[8][1] ),
    .A1(\rf.registers[9][1] ),
    .A2(\rf.registers[10][1] ),
    .A3(\rf.registers[11][1] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1136_));
 sky130_fd_sc_hd__mux4_2 _4381_ (.A0(\rf.registers[12][1] ),
    .A1(\rf.registers[13][1] ),
    .A2(\rf.registers[14][1] ),
    .A3(\rf.registers[15][1] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_2 _4382_ (.A0(_1136_),
    .A1(_1137_),
    .S(_1047_),
    .X(_1138_));
 sky130_fd_sc_hd__nand2_2 _4383_ (.A(_1038_),
    .B(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__mux4_2 _4384_ (.A0(\rf.registers[4][1] ),
    .A1(\rf.registers[5][1] ),
    .A2(\rf.registers[6][1] ),
    .A3(\rf.registers[7][1] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1140_));
 sky130_fd_sc_hd__mux4_2 _4385_ (.A0(\rf.registers[0][1] ),
    .A1(\rf.registers[1][1] ),
    .A2(\rf.registers[2][1] ),
    .A3(\rf.registers[3][1] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_2 _4386_ (.A0(_1140_),
    .A1(_1141_),
    .S(_1107_),
    .X(_1142_));
 sky130_fd_sc_hd__a21oi_2 _4387_ (.A1(_1088_),
    .A2(_1142_),
    .B1(A2[4]),
    .Y(_1143_));
 sky130_fd_sc_hd__a2bb2o_2 _4388_ (.A1_N(_1025_),
    .A2_N(_1135_),
    .B1(_1139_),
    .B2(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__buf_1 _4389_ (.A(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__buf_1 _4390_ (.A(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__buf_1 _4391_ (.A(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__buf_1 _4392_ (.A(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__buf_1 _4393_ (.A(A2[0]),
    .X(_1149_));
 sky130_fd_sc_hd__mux4_2 _4394_ (.A0(\rf.registers[20][0] ),
    .A1(\rf.registers[21][0] ),
    .A2(\rf.registers[22][0] ),
    .A3(\rf.registers[23][0] ),
    .S0(_1149_),
    .S1(_1061_),
    .X(_1150_));
 sky130_fd_sc_hd__mux4_2 _4395_ (.A0(\rf.registers[16][0] ),
    .A1(\rf.registers[17][0] ),
    .A2(\rf.registers[18][0] ),
    .A3(\rf.registers[19][0] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_2 _4396_ (.A0(_1150_),
    .A1(_1151_),
    .S(_1035_),
    .X(_1152_));
 sky130_fd_sc_hd__nand2_2 _4397_ (.A(_1088_),
    .B(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__mux4_2 _4398_ (.A0(\rf.registers[28][0] ),
    .A1(\rf.registers[29][0] ),
    .A2(\rf.registers[30][0] ),
    .A3(\rf.registers[31][0] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1154_));
 sky130_fd_sc_hd__mux4_2 _4399_ (.A0(\rf.registers[24][0] ),
    .A1(\rf.registers[25][0] ),
    .A2(\rf.registers[26][0] ),
    .A3(\rf.registers[27][0] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_2 _4400_ (.A0(_1154_),
    .A1(_1155_),
    .S(_1107_),
    .X(_1156_));
 sky130_fd_sc_hd__nand2_2 _4401_ (.A(_1038_),
    .B(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__mux4_2 _4402_ (.A0(\rf.registers[8][0] ),
    .A1(\rf.registers[9][0] ),
    .A2(\rf.registers[10][0] ),
    .A3(\rf.registers[11][0] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1158_));
 sky130_fd_sc_hd__mux4_2 _4403_ (.A0(\rf.registers[12][0] ),
    .A1(\rf.registers[13][0] ),
    .A2(\rf.registers[14][0] ),
    .A3(\rf.registers[15][0] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1159_));
 sky130_fd_sc_hd__mux2_2 _4404_ (.A0(_1158_),
    .A1(_1159_),
    .S(_1047_),
    .X(_1160_));
 sky130_fd_sc_hd__nand2_2 _4405_ (.A(_1038_),
    .B(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__mux4_2 _4406_ (.A0(\rf.registers[4][0] ),
    .A1(\rf.registers[5][0] ),
    .A2(\rf.registers[6][0] ),
    .A3(\rf.registers[7][0] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1162_));
 sky130_fd_sc_hd__mux4_2 _4407_ (.A0(\rf.registers[0][0] ),
    .A1(\rf.registers[1][0] ),
    .A2(\rf.registers[2][0] ),
    .A3(\rf.registers[3][0] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1163_));
 sky130_fd_sc_hd__mux2_2 _4408_ (.A0(_1162_),
    .A1(_1163_),
    .S(_1035_),
    .X(_1164_));
 sky130_fd_sc_hd__a21oi_2 _4409_ (.A1(_1088_),
    .A2(_1164_),
    .B1(A2[4]),
    .Y(_1165_));
 sky130_fd_sc_hd__a32o_2 _4410_ (.A1(_1057_),
    .A2(_1153_),
    .A3(_1157_),
    .B1(_1161_),
    .B2(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__buf_1 _4411_ (.A(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__buf_1 _4412_ (.A(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__buf_1 _4413_ (.A(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__buf_1 _4414_ (.A(_1057_),
    .X(_1170_));
 sky130_fd_sc_hd__buf_1 _4415_ (.A(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__buf_1 _4416_ (.A(_1072_),
    .X(_1172_));
 sky130_fd_sc_hd__buf_1 _4417_ (.A(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__buf_1 _4418_ (.A(_1073_),
    .X(_1174_));
 sky130_fd_sc_hd__buf_1 _4419_ (.A(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__mux4_2 _4420_ (.A0(\rf.registers[20][29] ),
    .A1(\rf.registers[21][29] ),
    .A2(\rf.registers[22][29] ),
    .A3(\rf.registers[23][29] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__mux4_2 _4421_ (.A0(\rf.registers[16][29] ),
    .A1(\rf.registers[17][29] ),
    .A2(\rf.registers[18][29] ),
    .A3(\rf.registers[19][29] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1177_));
 sky130_fd_sc_hd__buf_1 _4422_ (.A(_1036_),
    .X(_1178_));
 sky130_fd_sc_hd__mux2_2 _4423_ (.A0(_1176_),
    .A1(_1177_),
    .S(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__mux4_2 _4424_ (.A0(\rf.registers[28][29] ),
    .A1(\rf.registers[29][29] ),
    .A2(\rf.registers[30][29] ),
    .A3(\rf.registers[31][29] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1180_));
 sky130_fd_sc_hd__buf_1 _4425_ (.A(_1042_),
    .X(_1181_));
 sky130_fd_sc_hd__buf_1 _4426_ (.A(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__buf_1 _4427_ (.A(_1044_),
    .X(_1183_));
 sky130_fd_sc_hd__buf_1 _4428_ (.A(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__mux4_2 _4429_ (.A0(\rf.registers[24][29] ),
    .A1(\rf.registers[25][29] ),
    .A2(\rf.registers[26][29] ),
    .A3(\rf.registers[27][29] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__mux2_2 _4430_ (.A0(_1180_),
    .A1(_1185_),
    .S(_1178_),
    .X(_1186_));
 sky130_fd_sc_hd__buf_1 _4431_ (.A(_1071_),
    .X(_1187_));
 sky130_fd_sc_hd__mux2_2 _4432_ (.A0(_1179_),
    .A1(_1186_),
    .S(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__buf_1 _4433_ (.A(_1048_),
    .X(_1189_));
 sky130_fd_sc_hd__buf_1 _4434_ (.A(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__buf_1 _4435_ (.A(_1072_),
    .X(_1191_));
 sky130_fd_sc_hd__buf_1 _4436_ (.A(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__buf_1 _4437_ (.A(_1066_),
    .X(_1193_));
 sky130_fd_sc_hd__buf_1 _4438_ (.A(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__buf_1 _4439_ (.A(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__mux4_2 _4440_ (.A0(\rf.registers[12][29] ),
    .A1(\rf.registers[13][29] ),
    .A2(\rf.registers[14][29] ),
    .A3(\rf.registers[15][29] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__and2_2 _4441_ (.A(_1190_),
    .B(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__buf_1 _4442_ (.A(_1040_),
    .X(_1198_));
 sky130_fd_sc_hd__buf_1 _4443_ (.A(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__buf_1 _4444_ (.A(_1027_),
    .X(_1200_));
 sky130_fd_sc_hd__buf_1 _4445_ (.A(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__buf_1 _4446_ (.A(_1029_),
    .X(_1202_));
 sky130_fd_sc_hd__buf_1 _4447_ (.A(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__mux4_2 _4448_ (.A0(\rf.registers[8][29] ),
    .A1(\rf.registers[9][29] ),
    .A2(\rf.registers[10][29] ),
    .A3(\rf.registers[11][29] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__buf_1 _4449_ (.A(_1078_),
    .X(_1205_));
 sky130_fd_sc_hd__a21o_2 _4450_ (.A1(_1199_),
    .A2(_1204_),
    .B1(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__buf_1 _4451_ (.A(_1191_),
    .X(_1207_));
 sky130_fd_sc_hd__buf_1 _4452_ (.A(_1174_),
    .X(_1208_));
 sky130_fd_sc_hd__mux4_2 _4453_ (.A0(\rf.registers[4][29] ),
    .A1(\rf.registers[5][29] ),
    .A2(\rf.registers[6][29] ),
    .A3(\rf.registers[7][29] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__mux4_2 _4454_ (.A0(\rf.registers[0][29] ),
    .A1(\rf.registers[1][29] ),
    .A2(\rf.registers[2][29] ),
    .A3(\rf.registers[3][29] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1210_));
 sky130_fd_sc_hd__buf_1 _4455_ (.A(_1198_),
    .X(_1211_));
 sky130_fd_sc_hd__mux2_2 _4456_ (.A0(_1209_),
    .A1(_1210_),
    .S(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__buf_1 _4457_ (.A(_1038_),
    .X(_1213_));
 sky130_fd_sc_hd__buf_1 _4458_ (.A(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__buf_1 _4459_ (.A(_1025_),
    .X(_1215_));
 sky130_fd_sc_hd__o221a_2 _4460_ (.A1(_1197_),
    .A2(_1206_),
    .B1(_1212_),
    .B2(_1214_),
    .C1(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__a21oi_2 _4461_ (.A1(_1171_),
    .A2(_1188_),
    .B1(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__mux4_2 _4462_ (.A0(\rf.registers[20][28] ),
    .A1(\rf.registers[21][28] ),
    .A2(\rf.registers[22][28] ),
    .A3(\rf.registers[23][28] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1218_));
 sky130_fd_sc_hd__buf_1 _4463_ (.A(_1089_),
    .X(_1219_));
 sky130_fd_sc_hd__buf_1 _4464_ (.A(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__buf_1 _4465_ (.A(_1053_),
    .X(_1221_));
 sky130_fd_sc_hd__buf_1 _4466_ (.A(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__mux4_2 _4467_ (.A0(\rf.registers[16][28] ),
    .A1(\rf.registers[17][28] ),
    .A2(\rf.registers[18][28] ),
    .A3(\rf.registers[19][28] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_2 _4468_ (.A0(_1218_),
    .A1(_1223_),
    .S(_1178_),
    .X(_1224_));
 sky130_fd_sc_hd__mux4_2 _4469_ (.A0(\rf.registers[28][28] ),
    .A1(\rf.registers[29][28] ),
    .A2(\rf.registers[30][28] ),
    .A3(\rf.registers[31][28] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1225_));
 sky130_fd_sc_hd__mux4_2 _4470_ (.A0(\rf.registers[24][28] ),
    .A1(\rf.registers[25][28] ),
    .A2(\rf.registers[26][28] ),
    .A3(\rf.registers[27][28] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1226_));
 sky130_fd_sc_hd__mux2_2 _4471_ (.A0(_1225_),
    .A1(_1226_),
    .S(_1178_),
    .X(_1227_));
 sky130_fd_sc_hd__mux2_2 _4472_ (.A0(_1224_),
    .A1(_1227_),
    .S(_1187_),
    .X(_1228_));
 sky130_fd_sc_hd__mux4_2 _4473_ (.A0(\rf.registers[4][28] ),
    .A1(\rf.registers[5][28] ),
    .A2(\rf.registers[6][28] ),
    .A3(\rf.registers[7][28] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1229_));
 sky130_fd_sc_hd__and2_2 _4474_ (.A(_1189_),
    .B(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__mux4_2 _4475_ (.A0(\rf.registers[0][28] ),
    .A1(\rf.registers[1][28] ),
    .A2(\rf.registers[2][28] ),
    .A3(\rf.registers[3][28] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1231_));
 sky130_fd_sc_hd__a21o_2 _4476_ (.A1(_1199_),
    .A2(_1231_),
    .B1(_1213_),
    .X(_1232_));
 sky130_fd_sc_hd__mux4_2 _4477_ (.A0(\rf.registers[8][28] ),
    .A1(\rf.registers[9][28] ),
    .A2(\rf.registers[10][28] ),
    .A3(\rf.registers[11][28] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1233_));
 sky130_fd_sc_hd__mux4_2 _4478_ (.A0(\rf.registers[12][28] ),
    .A1(\rf.registers[13][28] ),
    .A2(\rf.registers[14][28] ),
    .A3(\rf.registers[15][28] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_2 _4479_ (.A0(_1233_),
    .A1(_1234_),
    .S(_1189_),
    .X(_1235_));
 sky130_fd_sc_hd__o221a_2 _4480_ (.A1(_1230_),
    .A2(_1232_),
    .B1(_1235_),
    .B2(_1205_),
    .C1(_1215_),
    .X(_1236_));
 sky130_fd_sc_hd__a21oi_2 _4481_ (.A1(_1171_),
    .A2(_1228_),
    .B1(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_2 _4482_ (.A(_1217_),
    .B(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__buf_1 _4483_ (.A(_1215_),
    .X(_1239_));
 sky130_fd_sc_hd__mux4_2 _4484_ (.A0(\rf.registers[20][20] ),
    .A1(\rf.registers[21][20] ),
    .A2(\rf.registers[22][20] ),
    .A3(\rf.registers[23][20] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1240_));
 sky130_fd_sc_hd__mux4_2 _4485_ (.A0(\rf.registers[16][20] ),
    .A1(\rf.registers[17][20] ),
    .A2(\rf.registers[18][20] ),
    .A3(\rf.registers[19][20] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_2 _4486_ (.A0(_1240_),
    .A1(_1241_),
    .S(_1211_),
    .X(_1242_));
 sky130_fd_sc_hd__mux4_2 _4487_ (.A0(\rf.registers[28][20] ),
    .A1(\rf.registers[29][20] ),
    .A2(\rf.registers[30][20] ),
    .A3(\rf.registers[31][20] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1243_));
 sky130_fd_sc_hd__mux4_2 _4488_ (.A0(\rf.registers[24][20] ),
    .A1(\rf.registers[25][20] ),
    .A2(\rf.registers[26][20] ),
    .A3(\rf.registers[27][20] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_2 _4489_ (.A0(_1243_),
    .A1(_1244_),
    .S(_1211_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_2 _4490_ (.A0(_1242_),
    .A1(_1245_),
    .S(_1187_),
    .X(_1246_));
 sky130_fd_sc_hd__mux4_2 _4491_ (.A0(\rf.registers[8][20] ),
    .A1(\rf.registers[9][20] ),
    .A2(\rf.registers[10][20] ),
    .A3(\rf.registers[11][20] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1247_));
 sky130_fd_sc_hd__or2_2 _4492_ (.A(_1190_),
    .B(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__mux4_2 _4493_ (.A0(\rf.registers[12][20] ),
    .A1(\rf.registers[13][20] ),
    .A2(\rf.registers[14][20] ),
    .A3(\rf.registers[15][20] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1249_));
 sky130_fd_sc_hd__o21a_2 _4494_ (.A1(_1199_),
    .A2(_1249_),
    .B1(_1213_),
    .X(_1250_));
 sky130_fd_sc_hd__mux4_2 _4495_ (.A0(\rf.registers[4][20] ),
    .A1(\rf.registers[5][20] ),
    .A2(\rf.registers[6][20] ),
    .A3(\rf.registers[7][20] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1251_));
 sky130_fd_sc_hd__mux4_2 _4496_ (.A0(\rf.registers[0][20] ),
    .A1(\rf.registers[1][20] ),
    .A2(\rf.registers[2][20] ),
    .A3(\rf.registers[3][20] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_2 _4497_ (.A0(_1251_),
    .A1(_1252_),
    .S(_1211_),
    .X(_1253_));
 sky130_fd_sc_hd__buf_1 _4498_ (.A(_1205_),
    .X(_1254_));
 sky130_fd_sc_hd__a221o_2 _4499_ (.A1(_1248_),
    .A2(_1250_),
    .B1(_1253_),
    .B2(_1254_),
    .C1(_1170_),
    .X(_1255_));
 sky130_fd_sc_hd__o21ai_2 _4500_ (.A1(_1239_),
    .A2(_1246_),
    .B1(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__mux4_2 _4501_ (.A0(\rf.registers[20][21] ),
    .A1(\rf.registers[21][21] ),
    .A2(\rf.registers[22][21] ),
    .A3(\rf.registers[23][21] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1257_));
 sky130_fd_sc_hd__mux4_2 _4502_ (.A0(\rf.registers[16][21] ),
    .A1(\rf.registers[17][21] ),
    .A2(\rf.registers[18][21] ),
    .A3(\rf.registers[19][21] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1258_));
 sky130_fd_sc_hd__buf_1 _4503_ (.A(_1036_),
    .X(_1259_));
 sky130_fd_sc_hd__mux2_2 _4504_ (.A0(_1257_),
    .A1(_1258_),
    .S(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__mux4_2 _4505_ (.A0(\rf.registers[28][21] ),
    .A1(\rf.registers[29][21] ),
    .A2(\rf.registers[30][21] ),
    .A3(\rf.registers[31][21] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1261_));
 sky130_fd_sc_hd__buf_1 _4506_ (.A(_1219_),
    .X(_1262_));
 sky130_fd_sc_hd__buf_1 _4507_ (.A(_1221_),
    .X(_1263_));
 sky130_fd_sc_hd__mux4_2 _4508_ (.A0(\rf.registers[24][21] ),
    .A1(\rf.registers[25][21] ),
    .A2(\rf.registers[26][21] ),
    .A3(\rf.registers[27][21] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_2 _4509_ (.A0(_1261_),
    .A1(_1264_),
    .S(_1259_),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_2 _4510_ (.A0(_1260_),
    .A1(_1265_),
    .S(_1187_),
    .X(_1266_));
 sky130_fd_sc_hd__buf_1 _4511_ (.A(_1200_),
    .X(_1267_));
 sky130_fd_sc_hd__buf_1 _4512_ (.A(_1202_),
    .X(_1268_));
 sky130_fd_sc_hd__mux4_2 _4513_ (.A0(\rf.registers[8][21] ),
    .A1(\rf.registers[9][21] ),
    .A2(\rf.registers[10][21] ),
    .A3(\rf.registers[11][21] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__mux4_2 _4514_ (.A0(\rf.registers[12][21] ),
    .A1(\rf.registers[13][21] ),
    .A2(\rf.registers[14][21] ),
    .A3(\rf.registers[15][21] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_2 _4515_ (.A0(_1269_),
    .A1(_1270_),
    .S(_1190_),
    .X(_1271_));
 sky130_fd_sc_hd__nand2_2 _4516_ (.A(_1214_),
    .B(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__mux4_2 _4517_ (.A0(\rf.registers[4][21] ),
    .A1(\rf.registers[5][21] ),
    .A2(\rf.registers[6][21] ),
    .A3(\rf.registers[7][21] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1273_));
 sky130_fd_sc_hd__mux4_2 _4518_ (.A0(\rf.registers[0][21] ),
    .A1(\rf.registers[1][21] ),
    .A2(\rf.registers[2][21] ),
    .A3(\rf.registers[3][21] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_2 _4519_ (.A0(_1273_),
    .A1(_1274_),
    .S(_1211_),
    .X(_1275_));
 sky130_fd_sc_hd__a21oi_2 _4520_ (.A1(_1254_),
    .A2(_1275_),
    .B1(_1171_),
    .Y(_1276_));
 sky130_fd_sc_hd__a2bb2o_2 _4521_ (.A1_N(_1239_),
    .A2_N(_1266_),
    .B1(_1272_),
    .B2(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__nand2_2 _4522_ (.A(_1256_),
    .B(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__buf_1 _4523_ (.A(_1073_),
    .X(_1279_));
 sky130_fd_sc_hd__mux4_2 _4524_ (.A0(\rf.registers[20][26] ),
    .A1(\rf.registers[21][26] ),
    .A2(\rf.registers[22][26] ),
    .A3(\rf.registers[23][26] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__mux4_2 _4525_ (.A0(\rf.registers[16][26] ),
    .A1(\rf.registers[17][26] ),
    .A2(\rf.registers[18][26] ),
    .A3(\rf.registers[19][26] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_2 _4526_ (.A0(_1280_),
    .A1(_1281_),
    .S(_1198_),
    .X(_1282_));
 sky130_fd_sc_hd__mux4_2 _4527_ (.A0(\rf.registers[28][26] ),
    .A1(\rf.registers[29][26] ),
    .A2(\rf.registers[30][26] ),
    .A3(\rf.registers[31][26] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1283_));
 sky130_fd_sc_hd__mux4_2 _4528_ (.A0(\rf.registers[24][26] ),
    .A1(\rf.registers[25][26] ),
    .A2(\rf.registers[26][26] ),
    .A3(\rf.registers[27][26] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1284_));
 sky130_fd_sc_hd__mux2_2 _4529_ (.A0(_1283_),
    .A1(_1284_),
    .S(_1198_),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_2 _4530_ (.A0(_1282_),
    .A1(_1285_),
    .S(_1071_),
    .X(_1286_));
 sky130_fd_sc_hd__buf_1 _4531_ (.A(_1048_),
    .X(_1287_));
 sky130_fd_sc_hd__mux4_2 _4532_ (.A0(\rf.registers[4][26] ),
    .A1(\rf.registers[5][26] ),
    .A2(\rf.registers[6][26] ),
    .A3(\rf.registers[7][26] ),
    .S0(_1191_),
    .S1(_1174_),
    .X(_1288_));
 sky130_fd_sc_hd__and2_2 _4533_ (.A(_1287_),
    .B(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__buf_1 _4534_ (.A(_1065_),
    .X(_1290_));
 sky130_fd_sc_hd__buf_1 _4535_ (.A(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__mux4_2 _4536_ (.A0(\rf.registers[0][26] ),
    .A1(\rf.registers[1][26] ),
    .A2(\rf.registers[2][26] ),
    .A3(\rf.registers[3][26] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1292_));
 sky130_fd_sc_hd__a21o_2 _4537_ (.A1(_1198_),
    .A2(_1292_),
    .B1(_1071_),
    .X(_1293_));
 sky130_fd_sc_hd__mux4_2 _4538_ (.A0(\rf.registers[8][26] ),
    .A1(\rf.registers[9][26] ),
    .A2(\rf.registers[10][26] ),
    .A3(\rf.registers[11][26] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1294_));
 sky130_fd_sc_hd__mux4_2 _4539_ (.A0(\rf.registers[12][26] ),
    .A1(\rf.registers[13][26] ),
    .A2(\rf.registers[14][26] ),
    .A3(\rf.registers[15][26] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_2 _4540_ (.A0(_1294_),
    .A1(_1295_),
    .S(_1287_),
    .X(_1296_));
 sky130_fd_sc_hd__o221a_2 _4541_ (.A1(_1289_),
    .A2(_1293_),
    .B1(_1296_),
    .B2(_1205_),
    .C1(_1025_),
    .X(_1297_));
 sky130_fd_sc_hd__a21o_2 _4542_ (.A1(_1170_),
    .A2(_1286_),
    .B1(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__inv_2 _4543_ (.A(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__mux4_2 _4544_ (.A0(\rf.registers[20][27] ),
    .A1(\rf.registers[21][27] ),
    .A2(\rf.registers[22][27] ),
    .A3(\rf.registers[23][27] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1300_));
 sky130_fd_sc_hd__mux4_2 _4545_ (.A0(\rf.registers[16][27] ),
    .A1(\rf.registers[17][27] ),
    .A2(\rf.registers[18][27] ),
    .A3(\rf.registers[19][27] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1301_));
 sky130_fd_sc_hd__mux2_2 _4546_ (.A0(_1300_),
    .A1(_1301_),
    .S(_1259_),
    .X(_1302_));
 sky130_fd_sc_hd__mux4_2 _4547_ (.A0(\rf.registers[28][27] ),
    .A1(\rf.registers[29][27] ),
    .A2(\rf.registers[30][27] ),
    .A3(\rf.registers[31][27] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1303_));
 sky130_fd_sc_hd__mux4_2 _4548_ (.A0(\rf.registers[24][27] ),
    .A1(\rf.registers[25][27] ),
    .A2(\rf.registers[26][27] ),
    .A3(\rf.registers[27][27] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1304_));
 sky130_fd_sc_hd__mux2_2 _4549_ (.A0(_1303_),
    .A1(_1304_),
    .S(_1259_),
    .X(_1305_));
 sky130_fd_sc_hd__mux2_2 _4550_ (.A0(_1302_),
    .A1(_1305_),
    .S(_1187_),
    .X(_1306_));
 sky130_fd_sc_hd__mux4_2 _4551_ (.A0(\rf.registers[12][27] ),
    .A1(\rf.registers[13][27] ),
    .A2(\rf.registers[14][27] ),
    .A3(\rf.registers[15][27] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1307_));
 sky130_fd_sc_hd__mux4_2 _4552_ (.A0(\rf.registers[8][27] ),
    .A1(\rf.registers[9][27] ),
    .A2(\rf.registers[10][27] ),
    .A3(\rf.registers[11][27] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_2 _4553_ (.A0(_1307_),
    .A1(_1308_),
    .S(_1199_),
    .X(_1309_));
 sky130_fd_sc_hd__nor2_2 _4554_ (.A(_1254_),
    .B(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__mux4_2 _4555_ (.A0(\rf.registers[4][27] ),
    .A1(\rf.registers[5][27] ),
    .A2(\rf.registers[6][27] ),
    .A3(\rf.registers[7][27] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1311_));
 sky130_fd_sc_hd__mux4_2 _4556_ (.A0(\rf.registers[0][27] ),
    .A1(\rf.registers[1][27] ),
    .A2(\rf.registers[2][27] ),
    .A3(\rf.registers[3][27] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1312_));
 sky130_fd_sc_hd__mux2_2 _4557_ (.A0(_1311_),
    .A1(_1312_),
    .S(_1199_),
    .X(_1313_));
 sky130_fd_sc_hd__o21ai_2 _4558_ (.A1(_1214_),
    .A2(_1313_),
    .B1(_1239_),
    .Y(_1314_));
 sky130_fd_sc_hd__o2bb2a_2 _4559_ (.A1_N(_1171_),
    .A2_N(_1306_),
    .B1(_1310_),
    .B2(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__nand2_2 _4560_ (.A(_1299_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__mux4_2 _4561_ (.A0(\rf.registers[20][31] ),
    .A1(\rf.registers[21][31] ),
    .A2(\rf.registers[22][31] ),
    .A3(\rf.registers[23][31] ),
    .S0(_1200_),
    .S1(_1202_),
    .X(_1317_));
 sky130_fd_sc_hd__mux4_2 _4562_ (.A0(\rf.registers[16][31] ),
    .A1(\rf.registers[17][31] ),
    .A2(\rf.registers[18][31] ),
    .A3(\rf.registers[19][31] ),
    .S0(_1200_),
    .S1(_1202_),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_2 _4563_ (.A0(_1317_),
    .A1(_1318_),
    .S(_1198_),
    .X(_1319_));
 sky130_fd_sc_hd__mux4_2 _4564_ (.A0(\rf.registers[28][31] ),
    .A1(\rf.registers[29][31] ),
    .A2(\rf.registers[30][31] ),
    .A3(\rf.registers[31][31] ),
    .S0(_1200_),
    .S1(_1202_),
    .X(_1320_));
 sky130_fd_sc_hd__mux4_2 _4565_ (.A0(\rf.registers[24][31] ),
    .A1(\rf.registers[25][31] ),
    .A2(\rf.registers[26][31] ),
    .A3(\rf.registers[27][31] ),
    .S0(_1200_),
    .S1(_1202_),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_2 _4566_ (.A0(_1320_),
    .A1(_1321_),
    .S(_1198_),
    .X(_1322_));
 sky130_fd_sc_hd__mux2_2 _4567_ (.A0(_1319_),
    .A1(_1322_),
    .S(_1213_),
    .X(_1323_));
 sky130_fd_sc_hd__buf_1 _4568_ (.A(_1027_),
    .X(_1324_));
 sky130_fd_sc_hd__buf_1 _4569_ (.A(_1029_),
    .X(_1325_));
 sky130_fd_sc_hd__mux4_2 _4570_ (.A0(\rf.registers[8][31] ),
    .A1(\rf.registers[9][31] ),
    .A2(\rf.registers[10][31] ),
    .A3(\rf.registers[11][31] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__and2_2 _4571_ (.A(_1178_),
    .B(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__mux4_2 _4572_ (.A0(\rf.registers[12][31] ),
    .A1(\rf.registers[13][31] ),
    .A2(\rf.registers[14][31] ),
    .A3(\rf.registers[15][31] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1328_));
 sky130_fd_sc_hd__a21o_2 _4573_ (.A1(_1189_),
    .A2(_1328_),
    .B1(_1078_),
    .X(_1329_));
 sky130_fd_sc_hd__mux4_2 _4574_ (.A0(\rf.registers[4][31] ),
    .A1(\rf.registers[5][31] ),
    .A2(\rf.registers[6][31] ),
    .A3(\rf.registers[7][31] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1330_));
 sky130_fd_sc_hd__mux4_2 _4575_ (.A0(\rf.registers[0][31] ),
    .A1(\rf.registers[1][31] ),
    .A2(\rf.registers[2][31] ),
    .A3(\rf.registers[3][31] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1331_));
 sky130_fd_sc_hd__mux2_2 _4576_ (.A0(_1330_),
    .A1(_1331_),
    .S(_1259_),
    .X(_1332_));
 sky130_fd_sc_hd__o221a_2 _4577_ (.A1(_1327_),
    .A2(_1329_),
    .B1(_1332_),
    .B2(_1187_),
    .C1(_1215_),
    .X(_1333_));
 sky130_fd_sc_hd__a21o_2 _4578_ (.A1(_1171_),
    .A2(_1323_),
    .B1(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__mux4_2 _4579_ (.A0(\rf.registers[24][30] ),
    .A1(\rf.registers[25][30] ),
    .A2(\rf.registers[26][30] ),
    .A3(\rf.registers[27][30] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1335_));
 sky130_fd_sc_hd__mux4_2 _4580_ (.A0(\rf.registers[28][30] ),
    .A1(\rf.registers[29][30] ),
    .A2(\rf.registers[30][30] ),
    .A3(\rf.registers[31][30] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1336_));
 sky130_fd_sc_hd__mux4_2 _4581_ (.A0(\rf.registers[16][30] ),
    .A1(\rf.registers[17][30] ),
    .A2(\rf.registers[18][30] ),
    .A3(\rf.registers[19][30] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1337_));
 sky130_fd_sc_hd__mux4_2 _4582_ (.A0(\rf.registers[20][30] ),
    .A1(\rf.registers[21][30] ),
    .A2(\rf.registers[22][30] ),
    .A3(\rf.registers[23][30] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1338_));
 sky130_fd_sc_hd__mux4_2 _4583_ (.A0(_1335_),
    .A1(_1336_),
    .A2(_1337_),
    .A3(_1338_),
    .S0(_1189_),
    .S1(_1205_),
    .X(_1339_));
 sky130_fd_sc_hd__mux4_2 _4584_ (.A0(\rf.registers[12][30] ),
    .A1(\rf.registers[13][30] ),
    .A2(\rf.registers[14][30] ),
    .A3(\rf.registers[15][30] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1340_));
 sky130_fd_sc_hd__and2_2 _4585_ (.A(_1189_),
    .B(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__mux4_2 _4586_ (.A0(\rf.registers[8][30] ),
    .A1(\rf.registers[9][30] ),
    .A2(\rf.registers[10][30] ),
    .A3(\rf.registers[11][30] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1342_));
 sky130_fd_sc_hd__a21o_2 _4587_ (.A1(_1211_),
    .A2(_1342_),
    .B1(_1078_),
    .X(_1343_));
 sky130_fd_sc_hd__mux4_2 _4588_ (.A0(\rf.registers[4][30] ),
    .A1(\rf.registers[5][30] ),
    .A2(\rf.registers[6][30] ),
    .A3(\rf.registers[7][30] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1344_));
 sky130_fd_sc_hd__mux4_2 _4589_ (.A0(\rf.registers[0][30] ),
    .A1(\rf.registers[1][30] ),
    .A2(\rf.registers[2][30] ),
    .A3(\rf.registers[3][30] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1345_));
 sky130_fd_sc_hd__mux2_2 _4590_ (.A0(_1344_),
    .A1(_1345_),
    .S(_1259_),
    .X(_1346_));
 sky130_fd_sc_hd__o221a_2 _4591_ (.A1(_1341_),
    .A2(_1343_),
    .B1(_1346_),
    .B2(_1187_),
    .C1(_1215_),
    .X(_1347_));
 sky130_fd_sc_hd__a21oi_2 _4592_ (.A1(_1171_),
    .A2(_1339_),
    .B1(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__or2b_2 _4593_ (.A(_1334_),
    .B_N(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__or4_2 _4594_ (.A(_1238_),
    .B(_1278_),
    .C(_1316_),
    .D(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__buf_1 _4595_ (.A(_1324_),
    .X(_1351_));
 sky130_fd_sc_hd__buf_1 _4596_ (.A(_1325_),
    .X(_1352_));
 sky130_fd_sc_hd__mux4_2 _4597_ (.A0(\rf.registers[20][25] ),
    .A1(\rf.registers[21][25] ),
    .A2(\rf.registers[22][25] ),
    .A3(\rf.registers[23][25] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__mux4_2 _4598_ (.A0(\rf.registers[16][25] ),
    .A1(\rf.registers[17][25] ),
    .A2(\rf.registers[18][25] ),
    .A3(\rf.registers[19][25] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1354_));
 sky130_fd_sc_hd__mux2_2 _4599_ (.A0(_1353_),
    .A1(_1354_),
    .S(_1199_),
    .X(_1355_));
 sky130_fd_sc_hd__mux4_2 _4600_ (.A0(\rf.registers[28][25] ),
    .A1(\rf.registers[29][25] ),
    .A2(\rf.registers[30][25] ),
    .A3(\rf.registers[31][25] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1356_));
 sky130_fd_sc_hd__mux4_2 _4601_ (.A0(\rf.registers[24][25] ),
    .A1(\rf.registers[25][25] ),
    .A2(\rf.registers[26][25] ),
    .A3(\rf.registers[27][25] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1357_));
 sky130_fd_sc_hd__mux2_2 _4602_ (.A0(_1356_),
    .A1(_1357_),
    .S(_1199_),
    .X(_1358_));
 sky130_fd_sc_hd__mux2_2 _4603_ (.A0(_1355_),
    .A1(_1358_),
    .S(_1214_),
    .X(_1359_));
 sky130_fd_sc_hd__buf_1 _4604_ (.A(_1351_),
    .X(_1360_));
 sky130_fd_sc_hd__buf_1 _4605_ (.A(_1352_),
    .X(_1361_));
 sky130_fd_sc_hd__mux4_2 _4606_ (.A0(\rf.registers[8][25] ),
    .A1(\rf.registers[9][25] ),
    .A2(\rf.registers[10][25] ),
    .A3(\rf.registers[11][25] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__mux4_2 _4607_ (.A0(\rf.registers[12][25] ),
    .A1(\rf.registers[13][25] ),
    .A2(\rf.registers[14][25] ),
    .A3(\rf.registers[15][25] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1363_));
 sky130_fd_sc_hd__mux2_2 _4608_ (.A0(_1362_),
    .A1(_1363_),
    .S(_1190_),
    .X(_1364_));
 sky130_fd_sc_hd__nor2_2 _4609_ (.A(_1254_),
    .B(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__mux4_2 _4610_ (.A0(\rf.registers[4][25] ),
    .A1(\rf.registers[5][25] ),
    .A2(\rf.registers[6][25] ),
    .A3(\rf.registers[7][25] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1366_));
 sky130_fd_sc_hd__mux4_2 _4611_ (.A0(\rf.registers[0][25] ),
    .A1(\rf.registers[1][25] ),
    .A2(\rf.registers[2][25] ),
    .A3(\rf.registers[3][25] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1367_));
 sky130_fd_sc_hd__mux2_2 _4612_ (.A0(_1366_),
    .A1(_1367_),
    .S(_1199_),
    .X(_1368_));
 sky130_fd_sc_hd__o21ai_2 _4613_ (.A1(_1214_),
    .A2(_1368_),
    .B1(_1239_),
    .Y(_1369_));
 sky130_fd_sc_hd__o2bb2a_2 _4614_ (.A1_N(_1171_),
    .A2_N(_1359_),
    .B1(_1365_),
    .B2(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__mux4_2 _4615_ (.A0(\rf.registers[24][24] ),
    .A1(\rf.registers[25][24] ),
    .A2(\rf.registers[26][24] ),
    .A3(\rf.registers[27][24] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1371_));
 sky130_fd_sc_hd__mux4_2 _4616_ (.A0(\rf.registers[28][24] ),
    .A1(\rf.registers[29][24] ),
    .A2(\rf.registers[30][24] ),
    .A3(\rf.registers[31][24] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1372_));
 sky130_fd_sc_hd__mux4_2 _4617_ (.A0(\rf.registers[16][24] ),
    .A1(\rf.registers[17][24] ),
    .A2(\rf.registers[18][24] ),
    .A3(\rf.registers[19][24] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1373_));
 sky130_fd_sc_hd__mux4_2 _4618_ (.A0(\rf.registers[20][24] ),
    .A1(\rf.registers[21][24] ),
    .A2(\rf.registers[22][24] ),
    .A3(\rf.registers[23][24] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1374_));
 sky130_fd_sc_hd__mux4_2 _4619_ (.A0(_1371_),
    .A1(_1372_),
    .A2(_1373_),
    .A3(_1374_),
    .S0(_1190_),
    .S1(_1254_),
    .X(_1375_));
 sky130_fd_sc_hd__mux4_2 _4620_ (.A0(\rf.registers[4][24] ),
    .A1(\rf.registers[5][24] ),
    .A2(\rf.registers[6][24] ),
    .A3(\rf.registers[7][24] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1376_));
 sky130_fd_sc_hd__mux4_2 _4621_ (.A0(\rf.registers[0][24] ),
    .A1(\rf.registers[1][24] ),
    .A2(\rf.registers[2][24] ),
    .A3(\rf.registers[3][24] ),
    .S0(_1360_),
    .S1(_1361_),
    .X(_1377_));
 sky130_fd_sc_hd__mux2_2 _4622_ (.A0(_1376_),
    .A1(_1377_),
    .S(_1199_),
    .X(_1378_));
 sky130_fd_sc_hd__nor2_2 _4623_ (.A(_1214_),
    .B(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__mux4_2 _4624_ (.A0(\rf.registers[8][24] ),
    .A1(\rf.registers[9][24] ),
    .A2(\rf.registers[10][24] ),
    .A3(\rf.registers[11][24] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1380_));
 sky130_fd_sc_hd__mux4_2 _4625_ (.A0(\rf.registers[12][24] ),
    .A1(\rf.registers[13][24] ),
    .A2(\rf.registers[14][24] ),
    .A3(\rf.registers[15][24] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1381_));
 sky130_fd_sc_hd__mux2_2 _4626_ (.A0(_1380_),
    .A1(_1381_),
    .S(_1190_),
    .X(_1382_));
 sky130_fd_sc_hd__o21ai_2 _4627_ (.A1(_1254_),
    .A2(_1382_),
    .B1(_1239_),
    .Y(_1383_));
 sky130_fd_sc_hd__o2bb2a_2 _4628_ (.A1_N(_1171_),
    .A2_N(_1375_),
    .B1(_1379_),
    .B2(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__nand2_2 _4629_ (.A(_1370_),
    .B(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__mux4_2 _4630_ (.A0(\rf.registers[24][6] ),
    .A1(\rf.registers[25][6] ),
    .A2(\rf.registers[26][6] ),
    .A3(\rf.registers[27][6] ),
    .S0(_1219_),
    .S1(_1221_),
    .X(_1386_));
 sky130_fd_sc_hd__mux4_2 _4631_ (.A0(\rf.registers[28][6] ),
    .A1(\rf.registers[29][6] ),
    .A2(\rf.registers[30][6] ),
    .A3(\rf.registers[31][6] ),
    .S0(_1219_),
    .S1(_1221_),
    .X(_1387_));
 sky130_fd_sc_hd__mux4_2 _4632_ (.A0(\rf.registers[16][6] ),
    .A1(\rf.registers[17][6] ),
    .A2(\rf.registers[18][6] ),
    .A3(\rf.registers[19][6] ),
    .S0(_1219_),
    .S1(_1221_),
    .X(_1388_));
 sky130_fd_sc_hd__mux4_2 _4633_ (.A0(\rf.registers[20][6] ),
    .A1(\rf.registers[21][6] ),
    .A2(\rf.registers[22][6] ),
    .A3(\rf.registers[23][6] ),
    .S0(_1219_),
    .S1(_1221_),
    .X(_1389_));
 sky130_fd_sc_hd__mux4_2 _4634_ (.A0(_1386_),
    .A1(_1387_),
    .A2(_1388_),
    .A3(_1389_),
    .S0(_1048_),
    .S1(_1088_),
    .X(_1390_));
 sky130_fd_sc_hd__mux4_2 _4635_ (.A0(\rf.registers[8][6] ),
    .A1(\rf.registers[9][6] ),
    .A2(\rf.registers[10][6] ),
    .A3(\rf.registers[11][6] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1391_));
 sky130_fd_sc_hd__or2_2 _4636_ (.A(_1048_),
    .B(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__mux4_2 _4637_ (.A0(\rf.registers[12][6] ),
    .A1(\rf.registers[13][6] ),
    .A2(\rf.registers[14][6] ),
    .A3(\rf.registers[15][6] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1393_));
 sky130_fd_sc_hd__o21a_2 _4638_ (.A1(_1036_),
    .A2(_1393_),
    .B1(_1037_),
    .X(_1394_));
 sky130_fd_sc_hd__mux4_2 _4639_ (.A0(\rf.registers[4][6] ),
    .A1(\rf.registers[5][6] ),
    .A2(\rf.registers[6][6] ),
    .A3(\rf.registers[7][6] ),
    .S0(_1072_),
    .S1(_1073_),
    .X(_1395_));
 sky130_fd_sc_hd__mux4_2 _4640_ (.A0(\rf.registers[0][6] ),
    .A1(\rf.registers[1][6] ),
    .A2(\rf.registers[2][6] ),
    .A3(\rf.registers[3][6] ),
    .S0(_1072_),
    .S1(_1073_),
    .X(_1396_));
 sky130_fd_sc_hd__mux2_2 _4641_ (.A0(_1395_),
    .A1(_1396_),
    .S(_1040_),
    .X(_1397_));
 sky130_fd_sc_hd__a221o_2 _4642_ (.A1(_1392_),
    .A2(_1394_),
    .B1(_1397_),
    .B2(_1078_),
    .C1(_1057_),
    .X(_1398_));
 sky130_fd_sc_hd__o21ai_2 _4643_ (.A1(_1025_),
    .A2(_1390_),
    .B1(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__mux4_2 _4644_ (.A0(\rf.registers[20][7] ),
    .A1(\rf.registers[21][7] ),
    .A2(\rf.registers[22][7] ),
    .A3(\rf.registers[23][7] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1400_));
 sky130_fd_sc_hd__mux4_2 _4645_ (.A0(\rf.registers[16][7] ),
    .A1(\rf.registers[17][7] ),
    .A2(\rf.registers[18][7] ),
    .A3(\rf.registers[19][7] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1401_));
 sky130_fd_sc_hd__mux2_2 _4646_ (.A0(_1400_),
    .A1(_1401_),
    .S(_1107_),
    .X(_1402_));
 sky130_fd_sc_hd__mux4_2 _4647_ (.A0(\rf.registers[28][7] ),
    .A1(\rf.registers[29][7] ),
    .A2(\rf.registers[30][7] ),
    .A3(\rf.registers[31][7] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1403_));
 sky130_fd_sc_hd__mux4_2 _4648_ (.A0(\rf.registers[24][7] ),
    .A1(\rf.registers[25][7] ),
    .A2(\rf.registers[26][7] ),
    .A3(\rf.registers[27][7] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_2 _4649_ (.A0(_1403_),
    .A1(_1404_),
    .S(_1107_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_2 _4650_ (.A0(_1402_),
    .A1(_1405_),
    .S(_1038_),
    .X(_1406_));
 sky130_fd_sc_hd__mux4_2 _4651_ (.A0(\rf.registers[12][7] ),
    .A1(\rf.registers[13][7] ),
    .A2(\rf.registers[14][7] ),
    .A3(\rf.registers[15][7] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1407_));
 sky130_fd_sc_hd__mux4_2 _4652_ (.A0(\rf.registers[8][7] ),
    .A1(\rf.registers[9][7] ),
    .A2(\rf.registers[10][7] ),
    .A3(\rf.registers[11][7] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1408_));
 sky130_fd_sc_hd__mux2_2 _4653_ (.A0(_1407_),
    .A1(_1408_),
    .S(_1040_),
    .X(_1409_));
 sky130_fd_sc_hd__nand2_2 _4654_ (.A(_1071_),
    .B(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__mux4_2 _4655_ (.A0(\rf.registers[4][7] ),
    .A1(\rf.registers[5][7] ),
    .A2(\rf.registers[6][7] ),
    .A3(\rf.registers[7][7] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1411_));
 sky130_fd_sc_hd__mux4_2 _4656_ (.A0(\rf.registers[0][7] ),
    .A1(\rf.registers[1][7] ),
    .A2(\rf.registers[2][7] ),
    .A3(\rf.registers[3][7] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_2 _4657_ (.A0(_1411_),
    .A1(_1412_),
    .S(_1040_),
    .X(_1413_));
 sky130_fd_sc_hd__a21oi_2 _4658_ (.A1(_1078_),
    .A2(_1413_),
    .B1(_1057_),
    .Y(_1414_));
 sky130_fd_sc_hd__a2bb2o_2 _4659_ (.A1_N(_1025_),
    .A2_N(_1406_),
    .B1(_1410_),
    .B2(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__nand2_2 _4660_ (.A(_1399_),
    .B(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__mux4_2 _4661_ (.A0(\rf.registers[24][23] ),
    .A1(\rf.registers[25][23] ),
    .A2(\rf.registers[26][23] ),
    .A3(\rf.registers[27][23] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1417_));
 sky130_fd_sc_hd__mux4_2 _4662_ (.A0(\rf.registers[28][23] ),
    .A1(\rf.registers[29][23] ),
    .A2(\rf.registers[30][23] ),
    .A3(\rf.registers[31][23] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1418_));
 sky130_fd_sc_hd__mux4_2 _4663_ (.A0(\rf.registers[16][23] ),
    .A1(\rf.registers[17][23] ),
    .A2(\rf.registers[18][23] ),
    .A3(\rf.registers[19][23] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1419_));
 sky130_fd_sc_hd__mux4_2 _4664_ (.A0(\rf.registers[20][23] ),
    .A1(\rf.registers[21][23] ),
    .A2(\rf.registers[22][23] ),
    .A3(\rf.registers[23][23] ),
    .S0(_1351_),
    .S1(_1352_),
    .X(_1420_));
 sky130_fd_sc_hd__mux4_2 _4665_ (.A0(_1417_),
    .A1(_1418_),
    .A2(_1419_),
    .A3(_1420_),
    .S0(_1190_),
    .S1(_1205_),
    .X(_1421_));
 sky130_fd_sc_hd__mux4_2 _4666_ (.A0(\rf.registers[8][23] ),
    .A1(\rf.registers[9][23] ),
    .A2(\rf.registers[10][23] ),
    .A3(\rf.registers[11][23] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1422_));
 sky130_fd_sc_hd__mux4_2 _4667_ (.A0(\rf.registers[12][23] ),
    .A1(\rf.registers[13][23] ),
    .A2(\rf.registers[14][23] ),
    .A3(\rf.registers[15][23] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_2 _4668_ (.A0(_1422_),
    .A1(_1423_),
    .S(_1190_),
    .X(_1424_));
 sky130_fd_sc_hd__nand2_2 _4669_ (.A(_1214_),
    .B(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__mux4_2 _4670_ (.A0(\rf.registers[4][23] ),
    .A1(\rf.registers[5][23] ),
    .A2(\rf.registers[6][23] ),
    .A3(\rf.registers[7][23] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1426_));
 sky130_fd_sc_hd__mux4_2 _4671_ (.A0(\rf.registers[0][23] ),
    .A1(\rf.registers[1][23] ),
    .A2(\rf.registers[2][23] ),
    .A3(\rf.registers[3][23] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1427_));
 sky130_fd_sc_hd__mux2_2 _4672_ (.A0(_1426_),
    .A1(_1427_),
    .S(_1211_),
    .X(_1428_));
 sky130_fd_sc_hd__a21oi_2 _4673_ (.A1(_1254_),
    .A2(_1428_),
    .B1(_1170_),
    .Y(_1429_));
 sky130_fd_sc_hd__a2bb2o_2 _4674_ (.A1_N(_1239_),
    .A2_N(_1421_),
    .B1(_1425_),
    .B2(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__mux4_2 _4675_ (.A0(\rf.registers[20][22] ),
    .A1(\rf.registers[21][22] ),
    .A2(\rf.registers[22][22] ),
    .A3(\rf.registers[23][22] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1431_));
 sky130_fd_sc_hd__mux4_2 _4676_ (.A0(\rf.registers[16][22] ),
    .A1(\rf.registers[17][22] ),
    .A2(\rf.registers[18][22] ),
    .A3(\rf.registers[19][22] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1432_));
 sky130_fd_sc_hd__mux2_2 _4677_ (.A0(_1431_),
    .A1(_1432_),
    .S(_1178_),
    .X(_1433_));
 sky130_fd_sc_hd__mux4_2 _4678_ (.A0(\rf.registers[28][22] ),
    .A1(\rf.registers[29][22] ),
    .A2(\rf.registers[30][22] ),
    .A3(\rf.registers[31][22] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1434_));
 sky130_fd_sc_hd__mux4_2 _4679_ (.A0(\rf.registers[24][22] ),
    .A1(\rf.registers[25][22] ),
    .A2(\rf.registers[26][22] ),
    .A3(\rf.registers[27][22] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1435_));
 sky130_fd_sc_hd__mux2_2 _4680_ (.A0(_1434_),
    .A1(_1435_),
    .S(_1178_),
    .X(_1436_));
 sky130_fd_sc_hd__mux2_2 _4681_ (.A0(_1433_),
    .A1(_1436_),
    .S(_1187_),
    .X(_1437_));
 sky130_fd_sc_hd__mux4_2 _4682_ (.A0(\rf.registers[8][22] ),
    .A1(\rf.registers[9][22] ),
    .A2(\rf.registers[10][22] ),
    .A3(\rf.registers[11][22] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1438_));
 sky130_fd_sc_hd__or2_2 _4683_ (.A(_1189_),
    .B(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__mux4_2 _4684_ (.A0(\rf.registers[12][22] ),
    .A1(\rf.registers[13][22] ),
    .A2(\rf.registers[14][22] ),
    .A3(\rf.registers[15][22] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1440_));
 sky130_fd_sc_hd__o21a_2 _4685_ (.A1(_1199_),
    .A2(_1440_),
    .B1(_1213_),
    .X(_1441_));
 sky130_fd_sc_hd__mux4_2 _4686_ (.A0(\rf.registers[4][22] ),
    .A1(\rf.registers[5][22] ),
    .A2(\rf.registers[6][22] ),
    .A3(\rf.registers[7][22] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1442_));
 sky130_fd_sc_hd__mux4_2 _4687_ (.A0(\rf.registers[0][22] ),
    .A1(\rf.registers[1][22] ),
    .A2(\rf.registers[2][22] ),
    .A3(\rf.registers[3][22] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_2 _4688_ (.A0(_1442_),
    .A1(_1443_),
    .S(_1211_),
    .X(_1444_));
 sky130_fd_sc_hd__a221o_2 _4689_ (.A1(_1439_),
    .A2(_1441_),
    .B1(_1444_),
    .B2(_1254_),
    .C1(_1170_),
    .X(_1445_));
 sky130_fd_sc_hd__o21ai_2 _4690_ (.A1(_1239_),
    .A2(_1437_),
    .B1(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__and2_2 _4691_ (.A(_1430_),
    .B(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__or2b_2 _4692_ (.A(_1416_),
    .B_N(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__mux4_2 _4693_ (.A0(\rf.registers[20][12] ),
    .A1(\rf.registers[21][12] ),
    .A2(\rf.registers[22][12] ),
    .A3(\rf.registers[23][12] ),
    .S0(_1219_),
    .S1(_1221_),
    .X(_1449_));
 sky130_fd_sc_hd__mux4_2 _4694_ (.A0(\rf.registers[16][12] ),
    .A1(\rf.registers[17][12] ),
    .A2(\rf.registers[18][12] ),
    .A3(\rf.registers[19][12] ),
    .S0(_1219_),
    .S1(_1221_),
    .X(_1450_));
 sky130_fd_sc_hd__mux2_2 _4695_ (.A0(_1449_),
    .A1(_1450_),
    .S(_1036_),
    .X(_1451_));
 sky130_fd_sc_hd__mux4_2 _4696_ (.A0(\rf.registers[28][12] ),
    .A1(\rf.registers[29][12] ),
    .A2(\rf.registers[30][12] ),
    .A3(\rf.registers[31][12] ),
    .S0(_1219_),
    .S1(_1221_),
    .X(_1452_));
 sky130_fd_sc_hd__mux4_2 _4697_ (.A0(\rf.registers[24][12] ),
    .A1(\rf.registers[25][12] ),
    .A2(\rf.registers[26][12] ),
    .A3(\rf.registers[27][12] ),
    .S0(_1219_),
    .S1(_1221_),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_2 _4698_ (.A0(_1452_),
    .A1(_1453_),
    .S(_1036_),
    .X(_1454_));
 sky130_fd_sc_hd__mux2_2 _4699_ (.A0(_1451_),
    .A1(_1454_),
    .S(_1071_),
    .X(_1455_));
 sky130_fd_sc_hd__mux4_2 _4700_ (.A0(\rf.registers[4][12] ),
    .A1(\rf.registers[5][12] ),
    .A2(\rf.registers[6][12] ),
    .A3(\rf.registers[7][12] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1456_));
 sky130_fd_sc_hd__or2_2 _4701_ (.A(_1198_),
    .B(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__mux4_2 _4702_ (.A0(\rf.registers[0][12] ),
    .A1(\rf.registers[1][12] ),
    .A2(\rf.registers[2][12] ),
    .A3(\rf.registers[3][12] ),
    .S0(_1191_),
    .S1(_1174_),
    .X(_1458_));
 sky130_fd_sc_hd__o21a_2 _4703_ (.A1(_1287_),
    .A2(_1458_),
    .B1(_1088_),
    .X(_1459_));
 sky130_fd_sc_hd__mux4_2 _4704_ (.A0(\rf.registers[8][12] ),
    .A1(\rf.registers[9][12] ),
    .A2(\rf.registers[10][12] ),
    .A3(\rf.registers[11][12] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1460_));
 sky130_fd_sc_hd__mux4_2 _4705_ (.A0(\rf.registers[12][12] ),
    .A1(\rf.registers[13][12] ),
    .A2(\rf.registers[14][12] ),
    .A3(\rf.registers[15][12] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_2 _4706_ (.A0(_1460_),
    .A1(_1461_),
    .S(_1048_),
    .X(_1462_));
 sky130_fd_sc_hd__a221o_2 _4707_ (.A1(_1457_),
    .A2(_1459_),
    .B1(_1462_),
    .B2(_1071_),
    .C1(_1057_),
    .X(_1463_));
 sky130_fd_sc_hd__o21ai_2 _4708_ (.A1(_1215_),
    .A2(_1455_),
    .B1(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__mux4_2 _4709_ (.A0(\rf.registers[20][13] ),
    .A1(\rf.registers[21][13] ),
    .A2(\rf.registers[22][13] ),
    .A3(\rf.registers[23][13] ),
    .S0(_1027_),
    .S1(_1029_),
    .X(_1465_));
 sky130_fd_sc_hd__mux4_2 _4710_ (.A0(\rf.registers[16][13] ),
    .A1(\rf.registers[17][13] ),
    .A2(\rf.registers[18][13] ),
    .A3(\rf.registers[19][13] ),
    .S0(_1027_),
    .S1(_1029_),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_2 _4711_ (.A0(_1465_),
    .A1(_1466_),
    .S(_1036_),
    .X(_1467_));
 sky130_fd_sc_hd__mux4_2 _4712_ (.A0(\rf.registers[28][13] ),
    .A1(\rf.registers[29][13] ),
    .A2(\rf.registers[30][13] ),
    .A3(\rf.registers[31][13] ),
    .S0(_1027_),
    .S1(_1029_),
    .X(_1468_));
 sky130_fd_sc_hd__mux4_2 _4713_ (.A0(\rf.registers[24][13] ),
    .A1(\rf.registers[25][13] ),
    .A2(\rf.registers[26][13] ),
    .A3(\rf.registers[27][13] ),
    .S0(_1027_),
    .S1(_1029_),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_2 _4714_ (.A0(_1468_),
    .A1(_1469_),
    .S(_1036_),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_2 _4715_ (.A0(_1467_),
    .A1(_1470_),
    .S(_1071_),
    .X(_1471_));
 sky130_fd_sc_hd__mux4_2 _4716_ (.A0(\rf.registers[8][13] ),
    .A1(\rf.registers[9][13] ),
    .A2(\rf.registers[10][13] ),
    .A3(\rf.registers[11][13] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1472_));
 sky130_fd_sc_hd__mux4_2 _4717_ (.A0(\rf.registers[12][13] ),
    .A1(\rf.registers[13][13] ),
    .A2(\rf.registers[14][13] ),
    .A3(\rf.registers[15][13] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_2 _4718_ (.A0(_1472_),
    .A1(_1473_),
    .S(_1287_),
    .X(_1474_));
 sky130_fd_sc_hd__nand2_2 _4719_ (.A(_1213_),
    .B(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__mux4_2 _4720_ (.A0(\rf.registers[4][13] ),
    .A1(\rf.registers[5][13] ),
    .A2(\rf.registers[6][13] ),
    .A3(\rf.registers[7][13] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1476_));
 sky130_fd_sc_hd__mux4_2 _4721_ (.A0(\rf.registers[0][13] ),
    .A1(\rf.registers[1][13] ),
    .A2(\rf.registers[2][13] ),
    .A3(\rf.registers[3][13] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_2 _4722_ (.A0(_1476_),
    .A1(_1477_),
    .S(_1198_),
    .X(_1478_));
 sky130_fd_sc_hd__a21oi_2 _4723_ (.A1(_1205_),
    .A2(_1478_),
    .B1(_1170_),
    .Y(_1479_));
 sky130_fd_sc_hd__a2bb2o_2 _4724_ (.A1_N(_1215_),
    .A2_N(_1471_),
    .B1(_1475_),
    .B2(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__mux4_2 _4725_ (.A0(\rf.registers[24][14] ),
    .A1(\rf.registers[25][14] ),
    .A2(\rf.registers[26][14] ),
    .A3(\rf.registers[27][14] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1481_));
 sky130_fd_sc_hd__mux4_2 _4726_ (.A0(\rf.registers[28][14] ),
    .A1(\rf.registers[29][14] ),
    .A2(\rf.registers[30][14] ),
    .A3(\rf.registers[31][14] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1482_));
 sky130_fd_sc_hd__mux4_2 _4727_ (.A0(\rf.registers[16][14] ),
    .A1(\rf.registers[17][14] ),
    .A2(\rf.registers[18][14] ),
    .A3(\rf.registers[19][14] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1483_));
 sky130_fd_sc_hd__mux4_2 _4728_ (.A0(\rf.registers[20][14] ),
    .A1(\rf.registers[21][14] ),
    .A2(\rf.registers[22][14] ),
    .A3(\rf.registers[23][14] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1484_));
 sky130_fd_sc_hd__mux4_2 _4729_ (.A0(_1481_),
    .A1(_1482_),
    .A2(_1483_),
    .A3(_1484_),
    .S0(_1189_),
    .S1(_1078_),
    .X(_1485_));
 sky130_fd_sc_hd__mux4_2 _4730_ (.A0(\rf.registers[4][14] ),
    .A1(\rf.registers[5][14] ),
    .A2(\rf.registers[6][14] ),
    .A3(\rf.registers[7][14] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1486_));
 sky130_fd_sc_hd__or2_2 _4731_ (.A(_1198_),
    .B(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__mux4_2 _4732_ (.A0(\rf.registers[0][14] ),
    .A1(\rf.registers[1][14] ),
    .A2(\rf.registers[2][14] ),
    .A3(\rf.registers[3][14] ),
    .S0(_1191_),
    .S1(_1174_),
    .X(_1488_));
 sky130_fd_sc_hd__o21a_2 _4733_ (.A1(_1287_),
    .A2(_1488_),
    .B1(_1078_),
    .X(_1489_));
 sky130_fd_sc_hd__mux4_2 _4734_ (.A0(\rf.registers[8][14] ),
    .A1(\rf.registers[9][14] ),
    .A2(\rf.registers[10][14] ),
    .A3(\rf.registers[11][14] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1490_));
 sky130_fd_sc_hd__mux4_2 _4735_ (.A0(\rf.registers[12][14] ),
    .A1(\rf.registers[13][14] ),
    .A2(\rf.registers[14][14] ),
    .A3(\rf.registers[15][14] ),
    .S0(_1172_),
    .S1(_1279_),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_2 _4736_ (.A0(_1490_),
    .A1(_1491_),
    .S(_1287_),
    .X(_1492_));
 sky130_fd_sc_hd__a221o_2 _4737_ (.A1(_1487_),
    .A2(_1489_),
    .B1(_1492_),
    .B2(_1213_),
    .C1(_1057_),
    .X(_1493_));
 sky130_fd_sc_hd__o21ai_2 _4738_ (.A1(_1215_),
    .A2(_1485_),
    .B1(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__and3_2 _4739_ (.A(_1464_),
    .B(_1480_),
    .C(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__mux4_2 _4740_ (.A0(\rf.registers[20][15] ),
    .A1(\rf.registers[21][15] ),
    .A2(\rf.registers[22][15] ),
    .A3(\rf.registers[23][15] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1496_));
 sky130_fd_sc_hd__mux4_2 _4741_ (.A0(\rf.registers[16][15] ),
    .A1(\rf.registers[17][15] ),
    .A2(\rf.registers[18][15] ),
    .A3(\rf.registers[19][15] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1497_));
 sky130_fd_sc_hd__mux2_2 _4742_ (.A0(_1496_),
    .A1(_1497_),
    .S(_1259_),
    .X(_1498_));
 sky130_fd_sc_hd__mux4_2 _4743_ (.A0(\rf.registers[28][15] ),
    .A1(\rf.registers[29][15] ),
    .A2(\rf.registers[30][15] ),
    .A3(\rf.registers[31][15] ),
    .S0(_1262_),
    .S1(_1263_),
    .X(_1499_));
 sky130_fd_sc_hd__mux4_2 _4744_ (.A0(\rf.registers[24][15] ),
    .A1(\rf.registers[25][15] ),
    .A2(\rf.registers[26][15] ),
    .A3(\rf.registers[27][15] ),
    .S0(_1324_),
    .S1(_1325_),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_2 _4745_ (.A0(_1499_),
    .A1(_1500_),
    .S(_1259_),
    .X(_1501_));
 sky130_fd_sc_hd__mux2_2 _4746_ (.A0(_1498_),
    .A1(_1501_),
    .S(_1187_),
    .X(_1502_));
 sky130_fd_sc_hd__mux4_2 _4747_ (.A0(\rf.registers[8][15] ),
    .A1(\rf.registers[9][15] ),
    .A2(\rf.registers[10][15] ),
    .A3(\rf.registers[11][15] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1503_));
 sky130_fd_sc_hd__mux4_2 _4748_ (.A0(\rf.registers[12][15] ),
    .A1(\rf.registers[13][15] ),
    .A2(\rf.registers[14][15] ),
    .A3(\rf.registers[15][15] ),
    .S0(_1201_),
    .S1(_1203_),
    .X(_1504_));
 sky130_fd_sc_hd__mux2_2 _4749_ (.A0(_1503_),
    .A1(_1504_),
    .S(_1190_),
    .X(_1505_));
 sky130_fd_sc_hd__nand2_2 _4750_ (.A(_1214_),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__mux4_2 _4751_ (.A0(\rf.registers[4][15] ),
    .A1(\rf.registers[5][15] ),
    .A2(\rf.registers[6][15] ),
    .A3(\rf.registers[7][15] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1507_));
 sky130_fd_sc_hd__mux4_2 _4752_ (.A0(\rf.registers[0][15] ),
    .A1(\rf.registers[1][15] ),
    .A2(\rf.registers[2][15] ),
    .A3(\rf.registers[3][15] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1508_));
 sky130_fd_sc_hd__mux2_2 _4753_ (.A0(_1507_),
    .A1(_1508_),
    .S(_1211_),
    .X(_1509_));
 sky130_fd_sc_hd__a21oi_2 _4754_ (.A1(_1254_),
    .A2(_1509_),
    .B1(_1170_),
    .Y(_1510_));
 sky130_fd_sc_hd__a2bb2o_2 _4755_ (.A1_N(_1239_),
    .A2_N(_1502_),
    .B1(_1506_),
    .B2(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__and2_2 _4756_ (.A(_1495_),
    .B(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__mux4_2 _4757_ (.A0(\rf.registers[20][8] ),
    .A1(\rf.registers[21][8] ),
    .A2(\rf.registers[22][8] ),
    .A3(\rf.registers[23][8] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1513_));
 sky130_fd_sc_hd__mux4_2 _4758_ (.A0(\rf.registers[16][8] ),
    .A1(\rf.registers[17][8] ),
    .A2(\rf.registers[18][8] ),
    .A3(\rf.registers[19][8] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1514_));
 sky130_fd_sc_hd__mux2_2 _4759_ (.A0(_1513_),
    .A1(_1514_),
    .S(_1035_),
    .X(_1515_));
 sky130_fd_sc_hd__mux4_2 _4760_ (.A0(\rf.registers[28][8] ),
    .A1(\rf.registers[29][8] ),
    .A2(\rf.registers[30][8] ),
    .A3(\rf.registers[31][8] ),
    .S0(_1026_),
    .S1(_1061_),
    .X(_1516_));
 sky130_fd_sc_hd__mux4_2 _4761_ (.A0(\rf.registers[24][8] ),
    .A1(\rf.registers[25][8] ),
    .A2(\rf.registers[26][8] ),
    .A3(\rf.registers[27][8] ),
    .S0(_1065_),
    .S1(_1066_),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_2 _4762_ (.A0(_1516_),
    .A1(_1517_),
    .S(_1035_),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_2 _4763_ (.A0(_1515_),
    .A1(_1518_),
    .S(_1037_),
    .X(_1519_));
 sky130_fd_sc_hd__mux4_2 _4764_ (.A0(\rf.registers[12][8] ),
    .A1(\rf.registers[13][8] ),
    .A2(\rf.registers[14][8] ),
    .A3(\rf.registers[15][8] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1520_));
 sky130_fd_sc_hd__or2_2 _4765_ (.A(_1107_),
    .B(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__mux4_2 _4766_ (.A0(\rf.registers[8][8] ),
    .A1(\rf.registers[9][8] ),
    .A2(\rf.registers[10][8] ),
    .A3(\rf.registers[11][8] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1522_));
 sky130_fd_sc_hd__o21a_2 _4767_ (.A1(_1047_),
    .A2(_1522_),
    .B1(_1037_),
    .X(_1523_));
 sky130_fd_sc_hd__mux4_2 _4768_ (.A0(\rf.registers[4][8] ),
    .A1(\rf.registers[5][8] ),
    .A2(\rf.registers[6][8] ),
    .A3(\rf.registers[7][8] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1524_));
 sky130_fd_sc_hd__mux4_2 _4769_ (.A0(\rf.registers[0][8] ),
    .A1(\rf.registers[1][8] ),
    .A2(\rf.registers[2][8] ),
    .A3(\rf.registers[3][8] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_2 _4770_ (.A0(_1524_),
    .A1(_1525_),
    .S(_1035_),
    .X(_1526_));
 sky130_fd_sc_hd__a221o_2 _4771_ (.A1(_1521_),
    .A2(_1523_),
    .B1(_1526_),
    .B2(_1050_),
    .C1(A2[4]),
    .X(_1527_));
 sky130_fd_sc_hd__o21a_2 _4772_ (.A1(_1025_),
    .A2(_1519_),
    .B1(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__mux4_2 _4773_ (.A0(\rf.registers[20][9] ),
    .A1(\rf.registers[21][9] ),
    .A2(\rf.registers[22][9] ),
    .A3(\rf.registers[23][9] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1529_));
 sky130_fd_sc_hd__mux4_2 _4774_ (.A0(\rf.registers[16][9] ),
    .A1(\rf.registers[17][9] ),
    .A2(\rf.registers[18][9] ),
    .A3(\rf.registers[19][9] ),
    .S0(_1072_),
    .S1(_1073_),
    .X(_1530_));
 sky130_fd_sc_hd__mux4_2 _4775_ (.A0(\rf.registers[28][9] ),
    .A1(\rf.registers[29][9] ),
    .A2(\rf.registers[30][9] ),
    .A3(\rf.registers[31][9] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1531_));
 sky130_fd_sc_hd__mux4_2 _4776_ (.A0(\rf.registers[24][9] ),
    .A1(\rf.registers[25][9] ),
    .A2(\rf.registers[26][9] ),
    .A3(\rf.registers[27][9] ),
    .S0(_1290_),
    .S1(_1193_),
    .X(_1532_));
 sky130_fd_sc_hd__mux4_2 _4777_ (.A0(_1529_),
    .A1(_1530_),
    .A2(_1531_),
    .A3(_1532_),
    .S0(_1040_),
    .S1(_1038_),
    .X(_1533_));
 sky130_fd_sc_hd__mux4_2 _4778_ (.A0(\rf.registers[8][9] ),
    .A1(\rf.registers[9][9] ),
    .A2(\rf.registers[10][9] ),
    .A3(\rf.registers[11][9] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1534_));
 sky130_fd_sc_hd__or2_2 _4779_ (.A(_1047_),
    .B(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__mux4_2 _4780_ (.A0(\rf.registers[12][9] ),
    .A1(\rf.registers[13][9] ),
    .A2(\rf.registers[14][9] ),
    .A3(\rf.registers[15][9] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1536_));
 sky130_fd_sc_hd__o21a_2 _4781_ (.A1(_1040_),
    .A2(_1536_),
    .B1(_1037_),
    .X(_1537_));
 sky130_fd_sc_hd__mux4_2 _4782_ (.A0(\rf.registers[4][9] ),
    .A1(\rf.registers[5][9] ),
    .A2(\rf.registers[6][9] ),
    .A3(\rf.registers[7][9] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1538_));
 sky130_fd_sc_hd__mux4_2 _4783_ (.A0(\rf.registers[0][9] ),
    .A1(\rf.registers[1][9] ),
    .A2(\rf.registers[2][9] ),
    .A3(\rf.registers[3][9] ),
    .S0(_1149_),
    .S1(_1028_),
    .X(_1539_));
 sky130_fd_sc_hd__mux2_2 _4784_ (.A0(_1538_),
    .A1(_1539_),
    .S(_1107_),
    .X(_1540_));
 sky130_fd_sc_hd__a221o_2 _4785_ (.A1(_1535_),
    .A2(_1537_),
    .B1(_1540_),
    .B2(_1088_),
    .C1(A2[4]),
    .X(_1541_));
 sky130_fd_sc_hd__o21ai_2 _4786_ (.A1(_1025_),
    .A2(_1533_),
    .B1(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__mux4_2 _4787_ (.A0(\rf.registers[20][10] ),
    .A1(\rf.registers[21][10] ),
    .A2(\rf.registers[22][10] ),
    .A3(\rf.registers[23][10] ),
    .S0(_1041_),
    .S1(_1043_),
    .X(_1543_));
 sky130_fd_sc_hd__mux4_2 _4788_ (.A0(\rf.registers[16][10] ),
    .A1(\rf.registers[17][10] ),
    .A2(\rf.registers[18][10] ),
    .A3(\rf.registers[19][10] ),
    .S0(_1041_),
    .S1(_1043_),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_2 _4789_ (.A0(_1543_),
    .A1(_1544_),
    .S(_1034_),
    .X(_1545_));
 sky130_fd_sc_hd__mux4_2 _4790_ (.A0(\rf.registers[28][10] ),
    .A1(\rf.registers[29][10] ),
    .A2(\rf.registers[30][10] ),
    .A3(\rf.registers[31][10] ),
    .S0(_1041_),
    .S1(_1043_),
    .X(_1546_));
 sky130_fd_sc_hd__mux4_2 _4791_ (.A0(\rf.registers[24][10] ),
    .A1(\rf.registers[25][10] ),
    .A2(\rf.registers[26][10] ),
    .A3(\rf.registers[27][10] ),
    .S0(_1041_),
    .S1(_1043_),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_2 _4792_ (.A0(_1546_),
    .A1(_1547_),
    .S(_1034_),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_2 _4793_ (.A0(_1545_),
    .A1(_1548_),
    .S(_1037_),
    .X(_1549_));
 sky130_fd_sc_hd__mux4_2 _4794_ (.A0(\rf.registers[8][10] ),
    .A1(\rf.registers[9][10] ),
    .A2(\rf.registers[10][10] ),
    .A3(\rf.registers[11][10] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1550_));
 sky130_fd_sc_hd__mux4_2 _4795_ (.A0(\rf.registers[12][10] ),
    .A1(\rf.registers[13][10] ),
    .A2(\rf.registers[14][10] ),
    .A3(\rf.registers[15][10] ),
    .S0(_1052_),
    .S1(_1090_),
    .X(_1551_));
 sky130_fd_sc_hd__mux2_2 _4796_ (.A0(_1550_),
    .A1(_1551_),
    .S(_1047_),
    .X(_1552_));
 sky130_fd_sc_hd__nand2_2 _4797_ (.A(_1038_),
    .B(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__mux4_2 _4798_ (.A0(\rf.registers[4][10] ),
    .A1(\rf.registers[5][10] ),
    .A2(\rf.registers[6][10] ),
    .A3(\rf.registers[7][10] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1554_));
 sky130_fd_sc_hd__mux4_2 _4799_ (.A0(\rf.registers[0][10] ),
    .A1(\rf.registers[1][10] ),
    .A2(\rf.registers[2][10] ),
    .A3(\rf.registers[3][10] ),
    .S0(_1104_),
    .S1(_1105_),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_2 _4800_ (.A0(_1554_),
    .A1(_1555_),
    .S(_1107_),
    .X(_1556_));
 sky130_fd_sc_hd__a21oi_2 _4801_ (.A1(_1088_),
    .A2(_1556_),
    .B1(A2[4]),
    .Y(_1557_));
 sky130_fd_sc_hd__a2bb2o_2 _4802_ (.A1_N(_1024_),
    .A2_N(_1549_),
    .B1(_1553_),
    .B2(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__mux4_2 _4803_ (.A0(\rf.registers[24][11] ),
    .A1(\rf.registers[25][11] ),
    .A2(\rf.registers[26][11] ),
    .A3(\rf.registers[27][11] ),
    .S0(_1072_),
    .S1(_1073_),
    .X(_1559_));
 sky130_fd_sc_hd__mux4_2 _4804_ (.A0(\rf.registers[28][11] ),
    .A1(\rf.registers[29][11] ),
    .A2(\rf.registers[30][11] ),
    .A3(\rf.registers[31][11] ),
    .S0(_1042_),
    .S1(_1044_),
    .X(_1560_));
 sky130_fd_sc_hd__mux4_2 _4805_ (.A0(\rf.registers[16][11] ),
    .A1(\rf.registers[17][11] ),
    .A2(\rf.registers[18][11] ),
    .A3(\rf.registers[19][11] ),
    .S0(_1072_),
    .S1(_1073_),
    .X(_1561_));
 sky130_fd_sc_hd__mux4_2 _4806_ (.A0(\rf.registers[20][11] ),
    .A1(\rf.registers[21][11] ),
    .A2(\rf.registers[22][11] ),
    .A3(\rf.registers[23][11] ),
    .S0(_1072_),
    .S1(_1073_),
    .X(_1562_));
 sky130_fd_sc_hd__mux4_2 _4807_ (.A0(_1559_),
    .A1(_1560_),
    .A2(_1561_),
    .A3(_1562_),
    .S0(_1048_),
    .S1(_1050_),
    .X(_1563_));
 sky130_fd_sc_hd__mux4_2 _4808_ (.A0(\rf.registers[8][11] ),
    .A1(\rf.registers[9][11] ),
    .A2(\rf.registers[10][11] ),
    .A3(\rf.registers[11][11] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1564_));
 sky130_fd_sc_hd__mux4_2 _4809_ (.A0(\rf.registers[12][11] ),
    .A1(\rf.registers[13][11] ),
    .A2(\rf.registers[14][11] ),
    .A3(\rf.registers[15][11] ),
    .S0(_1052_),
    .S1(_1053_),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_2 _4810_ (.A0(_1564_),
    .A1(_1565_),
    .S(_1048_),
    .X(_1566_));
 sky130_fd_sc_hd__nand2_2 _4811_ (.A(_1071_),
    .B(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__mux4_2 _4812_ (.A0(\rf.registers[4][11] ),
    .A1(\rf.registers[5][11] ),
    .A2(\rf.registers[6][11] ),
    .A3(\rf.registers[7][11] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1568_));
 sky130_fd_sc_hd__mux4_2 _4813_ (.A0(\rf.registers[0][11] ),
    .A1(\rf.registers[1][11] ),
    .A2(\rf.registers[2][11] ),
    .A3(\rf.registers[3][11] ),
    .S0(_1089_),
    .S1(_1090_),
    .X(_1569_));
 sky130_fd_sc_hd__mux2_2 _4814_ (.A0(_1568_),
    .A1(_1569_),
    .S(_1107_),
    .X(_1570_));
 sky130_fd_sc_hd__a21oi_2 _4815_ (.A1(_1088_),
    .A2(_1570_),
    .B1(A2[4]),
    .Y(_1571_));
 sky130_fd_sc_hd__a2bb2o_2 _4816_ (.A1_N(_1025_),
    .A2_N(_1563_),
    .B1(_1567_),
    .B2(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__and4b_2 _4817_ (.A_N(_1528_),
    .B(_1542_),
    .C(_1558_),
    .D(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__mux4_2 _4818_ (.A0(\rf.registers[24][16] ),
    .A1(\rf.registers[25][16] ),
    .A2(\rf.registers[26][16] ),
    .A3(\rf.registers[27][16] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1574_));
 sky130_fd_sc_hd__mux4_2 _4819_ (.A0(\rf.registers[28][16] ),
    .A1(\rf.registers[29][16] ),
    .A2(\rf.registers[30][16] ),
    .A3(\rf.registers[31][16] ),
    .S0(_1291_),
    .S1(_1174_),
    .X(_1575_));
 sky130_fd_sc_hd__mux4_2 _4820_ (.A0(\rf.registers[16][16] ),
    .A1(\rf.registers[17][16] ),
    .A2(\rf.registers[18][16] ),
    .A3(\rf.registers[19][16] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1576_));
 sky130_fd_sc_hd__mux4_2 _4821_ (.A0(\rf.registers[20][16] ),
    .A1(\rf.registers[21][16] ),
    .A2(\rf.registers[22][16] ),
    .A3(\rf.registers[23][16] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1577_));
 sky130_fd_sc_hd__mux4_2 _4822_ (.A0(_1574_),
    .A1(_1575_),
    .A2(_1576_),
    .A3(_1577_),
    .S0(_1287_),
    .S1(_1078_),
    .X(_1578_));
 sky130_fd_sc_hd__mux4_2 _4823_ (.A0(\rf.registers[8][16] ),
    .A1(\rf.registers[9][16] ),
    .A2(\rf.registers[10][16] ),
    .A3(\rf.registers[11][16] ),
    .S0(_1191_),
    .S1(_1174_),
    .X(_1579_));
 sky130_fd_sc_hd__mux4_2 _4824_ (.A0(\rf.registers[12][16] ),
    .A1(\rf.registers[13][16] ),
    .A2(\rf.registers[14][16] ),
    .A3(\rf.registers[15][16] ),
    .S0(_1191_),
    .S1(_1174_),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_2 _4825_ (.A0(_1579_),
    .A1(_1580_),
    .S(_1287_),
    .X(_1581_));
 sky130_fd_sc_hd__nand2_2 _4826_ (.A(_1213_),
    .B(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__mux4_2 _4827_ (.A0(\rf.registers[4][16] ),
    .A1(\rf.registers[5][16] ),
    .A2(\rf.registers[6][16] ),
    .A3(\rf.registers[7][16] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1583_));
 sky130_fd_sc_hd__mux4_2 _4828_ (.A0(\rf.registers[0][16] ),
    .A1(\rf.registers[1][16] ),
    .A2(\rf.registers[2][16] ),
    .A3(\rf.registers[3][16] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1584_));
 sky130_fd_sc_hd__mux2_2 _4829_ (.A0(_1583_),
    .A1(_1584_),
    .S(_1036_),
    .X(_1585_));
 sky130_fd_sc_hd__a21oi_2 _4830_ (.A1(_1205_),
    .A2(_1585_),
    .B1(_1170_),
    .Y(_1586_));
 sky130_fd_sc_hd__a2bb2o_2 _4831_ (.A1_N(_1215_),
    .A2_N(_1578_),
    .B1(_1582_),
    .B2(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__mux4_2 _4832_ (.A0(\rf.registers[24][17] ),
    .A1(\rf.registers[25][17] ),
    .A2(\rf.registers[26][17] ),
    .A3(\rf.registers[27][17] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1588_));
 sky130_fd_sc_hd__mux4_2 _4833_ (.A0(\rf.registers[28][17] ),
    .A1(\rf.registers[29][17] ),
    .A2(\rf.registers[30][17] ),
    .A3(\rf.registers[31][17] ),
    .S0(_1191_),
    .S1(_1174_),
    .X(_1589_));
 sky130_fd_sc_hd__mux4_2 _4834_ (.A0(\rf.registers[16][17] ),
    .A1(\rf.registers[17][17] ),
    .A2(\rf.registers[18][17] ),
    .A3(\rf.registers[19][17] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1590_));
 sky130_fd_sc_hd__mux4_2 _4835_ (.A0(\rf.registers[20][17] ),
    .A1(\rf.registers[21][17] ),
    .A2(\rf.registers[22][17] ),
    .A3(\rf.registers[23][17] ),
    .S0(_1291_),
    .S1(_1194_),
    .X(_1591_));
 sky130_fd_sc_hd__mux4_2 _4836_ (.A0(_1588_),
    .A1(_1589_),
    .A2(_1590_),
    .A3(_1591_),
    .S0(_1287_),
    .S1(_1078_),
    .X(_1592_));
 sky130_fd_sc_hd__mux4_2 _4837_ (.A0(\rf.registers[8][17] ),
    .A1(\rf.registers[9][17] ),
    .A2(\rf.registers[10][17] ),
    .A3(\rf.registers[11][17] ),
    .S0(_1191_),
    .S1(_1174_),
    .X(_1593_));
 sky130_fd_sc_hd__mux4_2 _4838_ (.A0(\rf.registers[12][17] ),
    .A1(\rf.registers[13][17] ),
    .A2(\rf.registers[14][17] ),
    .A3(\rf.registers[15][17] ),
    .S0(_1191_),
    .S1(_1279_),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_2 _4839_ (.A0(_1593_),
    .A1(_1594_),
    .S(_1287_),
    .X(_1595_));
 sky130_fd_sc_hd__nand2_2 _4840_ (.A(_1213_),
    .B(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__mux4_2 _4841_ (.A0(\rf.registers[4][17] ),
    .A1(\rf.registers[5][17] ),
    .A2(\rf.registers[6][17] ),
    .A3(\rf.registers[7][17] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1597_));
 sky130_fd_sc_hd__mux4_2 _4842_ (.A0(\rf.registers[0][17] ),
    .A1(\rf.registers[1][17] ),
    .A2(\rf.registers[2][17] ),
    .A3(\rf.registers[3][17] ),
    .S0(_1181_),
    .S1(_1183_),
    .X(_1598_));
 sky130_fd_sc_hd__mux2_2 _4843_ (.A0(_1597_),
    .A1(_1598_),
    .S(_1036_),
    .X(_1599_));
 sky130_fd_sc_hd__a21oi_2 _4844_ (.A1(_1205_),
    .A2(_1599_),
    .B1(_1057_),
    .Y(_1600_));
 sky130_fd_sc_hd__a2bb2o_2 _4845_ (.A1_N(_1215_),
    .A2_N(_1592_),
    .B1(_1596_),
    .B2(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__and2_2 _4846_ (.A(_1587_),
    .B(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__mux4_2 _4847_ (.A0(\rf.registers[20][19] ),
    .A1(\rf.registers[21][19] ),
    .A2(\rf.registers[22][19] ),
    .A3(\rf.registers[23][19] ),
    .S0(_1182_),
    .S1(_1184_),
    .X(_1603_));
 sky130_fd_sc_hd__mux4_2 _4848_ (.A0(\rf.registers[16][19] ),
    .A1(\rf.registers[17][19] ),
    .A2(\rf.registers[18][19] ),
    .A3(\rf.registers[19][19] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1604_));
 sky130_fd_sc_hd__mux2_2 _4849_ (.A0(_1603_),
    .A1(_1604_),
    .S(_1178_),
    .X(_1605_));
 sky130_fd_sc_hd__mux4_2 _4850_ (.A0(\rf.registers[28][19] ),
    .A1(\rf.registers[29][19] ),
    .A2(\rf.registers[30][19] ),
    .A3(\rf.registers[31][19] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1606_));
 sky130_fd_sc_hd__mux4_2 _4851_ (.A0(\rf.registers[24][19] ),
    .A1(\rf.registers[25][19] ),
    .A2(\rf.registers[26][19] ),
    .A3(\rf.registers[27][19] ),
    .S0(_1220_),
    .S1(_1222_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_2 _4852_ (.A0(_1606_),
    .A1(_1607_),
    .S(_1178_),
    .X(_1608_));
 sky130_fd_sc_hd__mux2_2 _4853_ (.A0(_1605_),
    .A1(_1608_),
    .S(_1187_),
    .X(_1609_));
 sky130_fd_sc_hd__mux4_2 _4854_ (.A0(\rf.registers[4][19] ),
    .A1(\rf.registers[5][19] ),
    .A2(\rf.registers[6][19] ),
    .A3(\rf.registers[7][19] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1610_));
 sky130_fd_sc_hd__or2_2 _4855_ (.A(_1211_),
    .B(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__mux4_2 _4856_ (.A0(\rf.registers[0][19] ),
    .A1(\rf.registers[1][19] ),
    .A2(\rf.registers[2][19] ),
    .A3(\rf.registers[3][19] ),
    .S0(_1207_),
    .S1(_1208_),
    .X(_1612_));
 sky130_fd_sc_hd__o21a_2 _4857_ (.A1(_1190_),
    .A2(_1612_),
    .B1(_1205_),
    .X(_1613_));
 sky130_fd_sc_hd__mux4_2 _4858_ (.A0(\rf.registers[8][19] ),
    .A1(\rf.registers[9][19] ),
    .A2(\rf.registers[10][19] ),
    .A3(\rf.registers[11][19] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1614_));
 sky130_fd_sc_hd__mux4_2 _4859_ (.A0(\rf.registers[12][19] ),
    .A1(\rf.registers[13][19] ),
    .A2(\rf.registers[14][19] ),
    .A3(\rf.registers[15][19] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1615_));
 sky130_fd_sc_hd__mux2_2 _4860_ (.A0(_1614_),
    .A1(_1615_),
    .S(_1189_),
    .X(_1616_));
 sky130_fd_sc_hd__a221o_2 _4861_ (.A1(_1611_),
    .A2(_1613_),
    .B1(_1616_),
    .B2(_1214_),
    .C1(_1170_),
    .X(_1617_));
 sky130_fd_sc_hd__o21ai_2 _4862_ (.A1(_1239_),
    .A2(_1609_),
    .B1(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__mux4_2 _4863_ (.A0(\rf.registers[20][18] ),
    .A1(\rf.registers[21][18] ),
    .A2(\rf.registers[22][18] ),
    .A3(\rf.registers[23][18] ),
    .S0(_1200_),
    .S1(_1202_),
    .X(_1619_));
 sky130_fd_sc_hd__mux4_2 _4864_ (.A0(\rf.registers[16][18] ),
    .A1(\rf.registers[17][18] ),
    .A2(\rf.registers[18][18] ),
    .A3(\rf.registers[19][18] ),
    .S0(_1200_),
    .S1(_1202_),
    .X(_1620_));
 sky130_fd_sc_hd__mux2_2 _4865_ (.A0(_1619_),
    .A1(_1620_),
    .S(_1259_),
    .X(_1621_));
 sky130_fd_sc_hd__mux4_2 _4866_ (.A0(\rf.registers[28][18] ),
    .A1(\rf.registers[29][18] ),
    .A2(\rf.registers[30][18] ),
    .A3(\rf.registers[31][18] ),
    .S0(_1200_),
    .S1(_1202_),
    .X(_1622_));
 sky130_fd_sc_hd__mux4_2 _4867_ (.A0(\rf.registers[24][18] ),
    .A1(\rf.registers[25][18] ),
    .A2(\rf.registers[26][18] ),
    .A3(\rf.registers[27][18] ),
    .S0(_1200_),
    .S1(_1202_),
    .X(_1623_));
 sky130_fd_sc_hd__mux2_2 _4868_ (.A0(_1622_),
    .A1(_1623_),
    .S(_1259_),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_2 _4869_ (.A0(_1621_),
    .A1(_1624_),
    .S(_1213_),
    .X(_1625_));
 sky130_fd_sc_hd__mux4_2 _4870_ (.A0(\rf.registers[8][18] ),
    .A1(\rf.registers[9][18] ),
    .A2(\rf.registers[10][18] ),
    .A3(\rf.registers[11][18] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1626_));
 sky130_fd_sc_hd__mux4_2 _4871_ (.A0(\rf.registers[12][18] ),
    .A1(\rf.registers[13][18] ),
    .A2(\rf.registers[14][18] ),
    .A3(\rf.registers[15][18] ),
    .S0(_1192_),
    .S1(_1195_),
    .X(_1627_));
 sky130_fd_sc_hd__mux2_2 _4872_ (.A0(_1626_),
    .A1(_1627_),
    .S(_1189_),
    .X(_1628_));
 sky130_fd_sc_hd__nand2_2 _4873_ (.A(_1214_),
    .B(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__mux4_2 _4874_ (.A0(\rf.registers[4][18] ),
    .A1(\rf.registers[5][18] ),
    .A2(\rf.registers[6][18] ),
    .A3(\rf.registers[7][18] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1630_));
 sky130_fd_sc_hd__mux4_2 _4875_ (.A0(\rf.registers[0][18] ),
    .A1(\rf.registers[1][18] ),
    .A2(\rf.registers[2][18] ),
    .A3(\rf.registers[3][18] ),
    .S0(_1173_),
    .S1(_1175_),
    .X(_1631_));
 sky130_fd_sc_hd__mux2_2 _4876_ (.A0(_1630_),
    .A1(_1631_),
    .S(_1178_),
    .X(_1632_));
 sky130_fd_sc_hd__a21oi_2 _4877_ (.A1(_1254_),
    .A2(_1632_),
    .B1(_1170_),
    .Y(_1633_));
 sky130_fd_sc_hd__a2bb2o_2 _4878_ (.A1_N(_1239_),
    .A2_N(_1625_),
    .B1(_1629_),
    .B2(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__and3_2 _4879_ (.A(_1602_),
    .B(_1618_),
    .C(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__and3_2 _4880_ (.A(_1512_),
    .B(_1573_),
    .C(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__or4b_2 _4881_ (.A(_1350_),
    .B(_1385_),
    .C(_1448_),
    .D_N(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__buf_1 _4882_ (.A(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__buf_1 _4883_ (.A(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__inv_2 _4884_ (.A(A1[4]),
    .Y(_1640_));
 sky130_fd_sc_hd__buf_1 _4885_ (.A(A1[0]),
    .X(_1641_));
 sky130_fd_sc_hd__buf_1 _4886_ (.A(A1[1]),
    .X(_1642_));
 sky130_fd_sc_hd__mux4_2 _4887_ (.A0(\rf.registers[20][0] ),
    .A1(\rf.registers[21][0] ),
    .A2(\rf.registers[22][0] ),
    .A3(\rf.registers[23][0] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__mux4_2 _4888_ (.A0(\rf.registers[16][0] ),
    .A1(\rf.registers[17][0] ),
    .A2(\rf.registers[18][0] ),
    .A3(\rf.registers[19][0] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_1644_));
 sky130_fd_sc_hd__inv_2 _4889_ (.A(A1[2]),
    .Y(_1645_));
 sky130_fd_sc_hd__mux2_2 _4890_ (.A0(_1643_),
    .A1(_1644_),
    .S(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__mux4_2 _4891_ (.A0(\rf.registers[28][0] ),
    .A1(\rf.registers[29][0] ),
    .A2(\rf.registers[30][0] ),
    .A3(\rf.registers[31][0] ),
    .S0(A1[0]),
    .S1(A1[1]),
    .X(_1647_));
 sky130_fd_sc_hd__mux4_2 _4892_ (.A0(\rf.registers[24][0] ),
    .A1(\rf.registers[25][0] ),
    .A2(\rf.registers[26][0] ),
    .A3(\rf.registers[27][0] ),
    .S0(A1[0]),
    .S1(A1[1]),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_2 _4893_ (.A0(_1647_),
    .A1(_1648_),
    .S(_1645_),
    .X(_1649_));
 sky130_fd_sc_hd__mux2_2 _4894_ (.A0(_1646_),
    .A1(_1649_),
    .S(A1[3]),
    .X(_1650_));
 sky130_fd_sc_hd__mux4_2 _4895_ (.A0(\rf.registers[8][0] ),
    .A1(\rf.registers[9][0] ),
    .A2(\rf.registers[10][0] ),
    .A3(\rf.registers[11][0] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_1651_));
 sky130_fd_sc_hd__mux4_2 _4896_ (.A0(\rf.registers[12][0] ),
    .A1(\rf.registers[13][0] ),
    .A2(\rf.registers[14][0] ),
    .A3(\rf.registers[15][0] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_1652_));
 sky130_fd_sc_hd__mux2_2 _4897_ (.A0(_1651_),
    .A1(_1652_),
    .S(A1[2]),
    .X(_1653_));
 sky130_fd_sc_hd__nand2_2 _4898_ (.A(A1[3]),
    .B(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__inv_2 _4899_ (.A(A1[3]),
    .Y(_1655_));
 sky130_fd_sc_hd__mux4_2 _4900_ (.A0(\rf.registers[4][0] ),
    .A1(\rf.registers[5][0] ),
    .A2(\rf.registers[6][0] ),
    .A3(\rf.registers[7][0] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_1656_));
 sky130_fd_sc_hd__mux4_2 _4901_ (.A0(\rf.registers[0][0] ),
    .A1(\rf.registers[1][0] ),
    .A2(\rf.registers[2][0] ),
    .A3(\rf.registers[3][0] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_1657_));
 sky130_fd_sc_hd__mux2_2 _4902_ (.A0(_1656_),
    .A1(_1657_),
    .S(_1645_),
    .X(_1658_));
 sky130_fd_sc_hd__a21oi_2 _4903_ (.A1(_1655_),
    .A2(_1658_),
    .B1(A1[4]),
    .Y(_1659_));
 sky130_fd_sc_hd__a2bb2o_2 _4904_ (.A1_N(_1640_),
    .A2_N(_1650_),
    .B1(_1654_),
    .B2(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__nor2_2 _4905_ (.A(_1639_),
    .B(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__and2_2 _4906_ (.A(_1169_),
    .B(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__nand2_2 _4907_ (.A(_1148_),
    .B(_1662_),
    .Y(_1663_));
 sky130_fd_sc_hd__inv_2 _4908_ (.A(opcode[0]),
    .Y(_1664_));
 sky130_fd_sc_hd__or3_2 _4909_ (.A(_1664_),
    .B(_1060_),
    .C(_1084_),
    .X(_1665_));
 sky130_fd_sc_hd__buf_1 _4910_ (.A(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__a32oi_2 _4911_ (.A1(_1171_),
    .A2(_1153_),
    .A3(_1157_),
    .B1(_1161_),
    .B2(_1165_),
    .Y(_1667_));
 sky130_fd_sc_hd__buf_1 _4912_ (.A(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__buf_1 _4913_ (.A(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__buf_1 _4914_ (.A(_1640_),
    .X(_1670_));
 sky130_fd_sc_hd__buf_1 _4915_ (.A(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__buf_1 _4916_ (.A(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__buf_1 _4917_ (.A(_1641_),
    .X(_1673_));
 sky130_fd_sc_hd__buf_1 _4918_ (.A(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__buf_1 _4919_ (.A(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__buf_1 _4920_ (.A(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__buf_1 _4921_ (.A(A1[1]),
    .X(_1677_));
 sky130_fd_sc_hd__buf_1 _4922_ (.A(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__buf_1 _4923_ (.A(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__buf_1 _4924_ (.A(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__buf_1 _4925_ (.A(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__mux4_2 _4926_ (.A0(\rf.registers[20][23] ),
    .A1(\rf.registers[21][23] ),
    .A2(\rf.registers[22][23] ),
    .A3(\rf.registers[23][23] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__mux4_2 _4927_ (.A0(\rf.registers[16][23] ),
    .A1(\rf.registers[17][23] ),
    .A2(\rf.registers[18][23] ),
    .A3(\rf.registers[19][23] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1683_));
 sky130_fd_sc_hd__buf_1 _4928_ (.A(_1645_),
    .X(_1684_));
 sky130_fd_sc_hd__buf_1 _4929_ (.A(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__buf_1 _4930_ (.A(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__mux2_2 _4931_ (.A0(_1682_),
    .A1(_1683_),
    .S(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__mux4_2 _4932_ (.A0(\rf.registers[28][23] ),
    .A1(\rf.registers[29][23] ),
    .A2(\rf.registers[30][23] ),
    .A3(\rf.registers[31][23] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1688_));
 sky130_fd_sc_hd__buf_1 _4933_ (.A(_1675_),
    .X(_1689_));
 sky130_fd_sc_hd__buf_1 _4934_ (.A(_1642_),
    .X(_1690_));
 sky130_fd_sc_hd__buf_1 _4935_ (.A(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__buf_1 _4936_ (.A(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__buf_1 _4937_ (.A(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__mux4_2 _4938_ (.A0(\rf.registers[24][23] ),
    .A1(\rf.registers[25][23] ),
    .A2(\rf.registers[26][23] ),
    .A3(\rf.registers[27][23] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__mux2_2 _4939_ (.A0(_1688_),
    .A1(_1694_),
    .S(_1686_),
    .X(_1695_));
 sky130_fd_sc_hd__buf_1 _4940_ (.A(A1[3]),
    .X(_1696_));
 sky130_fd_sc_hd__buf_1 _4941_ (.A(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__mux2_2 _4942_ (.A0(_1687_),
    .A1(_1695_),
    .S(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__buf_1 _4943_ (.A(_1696_),
    .X(_1699_));
 sky130_fd_sc_hd__buf_1 _4944_ (.A(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__buf_1 _4945_ (.A(A1[0]),
    .X(_1701_));
 sky130_fd_sc_hd__buf_1 _4946_ (.A(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__buf_1 _4947_ (.A(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__buf_1 _4948_ (.A(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__buf_1 _4949_ (.A(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__buf_1 _4950_ (.A(_1678_),
    .X(_1706_));
 sky130_fd_sc_hd__buf_1 _4951_ (.A(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__buf_1 _4952_ (.A(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__mux4_2 _4953_ (.A0(\rf.registers[8][23] ),
    .A1(\rf.registers[9][23] ),
    .A2(\rf.registers[10][23] ),
    .A3(\rf.registers[11][23] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__mux4_2 _4954_ (.A0(\rf.registers[12][23] ),
    .A1(\rf.registers[13][23] ),
    .A2(\rf.registers[14][23] ),
    .A3(\rf.registers[15][23] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1710_));
 sky130_fd_sc_hd__buf_1 _4955_ (.A(A1[2]),
    .X(_1711_));
 sky130_fd_sc_hd__buf_1 _4956_ (.A(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__buf_1 _4957_ (.A(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__mux2_2 _4958_ (.A0(_1709_),
    .A1(_1710_),
    .S(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__nand2_2 _4959_ (.A(_1700_),
    .B(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__buf_1 _4960_ (.A(_1655_),
    .X(_1716_));
 sky130_fd_sc_hd__buf_1 _4961_ (.A(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__buf_1 _4962_ (.A(_1702_),
    .X(_1718_));
 sky130_fd_sc_hd__buf_1 _4963_ (.A(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__buf_1 _4964_ (.A(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__buf_1 _4965_ (.A(_1678_),
    .X(_1721_));
 sky130_fd_sc_hd__buf_1 _4966_ (.A(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__buf_1 _4967_ (.A(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__mux4_2 _4968_ (.A0(\rf.registers[4][23] ),
    .A1(\rf.registers[5][23] ),
    .A2(\rf.registers[6][23] ),
    .A3(\rf.registers[7][23] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__mux4_2 _4969_ (.A0(\rf.registers[0][23] ),
    .A1(\rf.registers[1][23] ),
    .A2(\rf.registers[2][23] ),
    .A3(\rf.registers[3][23] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1725_));
 sky130_fd_sc_hd__buf_1 _4970_ (.A(_1685_),
    .X(_1726_));
 sky130_fd_sc_hd__mux2_2 _4971_ (.A0(_1724_),
    .A1(_1725_),
    .S(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__buf_1 _4972_ (.A(A1[4]),
    .X(_1728_));
 sky130_fd_sc_hd__buf_1 _4973_ (.A(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__a21oi_2 _4974_ (.A1(_1717_),
    .A2(_1727_),
    .B1(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__a2bb2o_2 _4975_ (.A1_N(_1672_),
    .A2_N(_1698_),
    .B1(_1715_),
    .B2(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__or2_2 _4976_ (.A(_1639_),
    .B(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__buf_1 _4977_ (.A(_1702_),
    .X(_1733_));
 sky130_fd_sc_hd__buf_1 _4978_ (.A(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__buf_1 _4979_ (.A(_1721_),
    .X(_1735_));
 sky130_fd_sc_hd__mux4_2 _4980_ (.A0(\rf.registers[20][22] ),
    .A1(\rf.registers[21][22] ),
    .A2(\rf.registers[22][22] ),
    .A3(\rf.registers[23][22] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__mux4_2 _4981_ (.A0(\rf.registers[16][22] ),
    .A1(\rf.registers[17][22] ),
    .A2(\rf.registers[18][22] ),
    .A3(\rf.registers[19][22] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_1737_));
 sky130_fd_sc_hd__buf_1 _4982_ (.A(_1684_),
    .X(_1738_));
 sky130_fd_sc_hd__buf_1 _4983_ (.A(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__mux2_2 _4984_ (.A0(_1736_),
    .A1(_1737_),
    .S(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__mux4_2 _4985_ (.A0(\rf.registers[28][22] ),
    .A1(\rf.registers[29][22] ),
    .A2(\rf.registers[30][22] ),
    .A3(\rf.registers[31][22] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_1741_));
 sky130_fd_sc_hd__mux4_2 _4986_ (.A0(\rf.registers[24][22] ),
    .A1(\rf.registers[25][22] ),
    .A2(\rf.registers[26][22] ),
    .A3(\rf.registers[27][22] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_1742_));
 sky130_fd_sc_hd__mux2_2 _4987_ (.A0(_1741_),
    .A1(_1742_),
    .S(_1739_),
    .X(_1743_));
 sky130_fd_sc_hd__mux2_2 _4988_ (.A0(_1740_),
    .A1(_1743_),
    .S(_1697_),
    .X(_1744_));
 sky130_fd_sc_hd__buf_1 _4989_ (.A(_1686_),
    .X(_1745_));
 sky130_fd_sc_hd__mux4_2 _4990_ (.A0(\rf.registers[12][22] ),
    .A1(\rf.registers[13][22] ),
    .A2(\rf.registers[14][22] ),
    .A3(\rf.registers[15][22] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1746_));
 sky130_fd_sc_hd__mux4_2 _4991_ (.A0(\rf.registers[8][22] ),
    .A1(\rf.registers[9][22] ),
    .A2(\rf.registers[10][22] ),
    .A3(\rf.registers[11][22] ),
    .S0(_1704_),
    .S1(_1707_),
    .X(_1747_));
 sky130_fd_sc_hd__or2_2 _4992_ (.A(_1712_),
    .B(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__o211a_2 _4993_ (.A1(_1745_),
    .A2(_1746_),
    .B1(_1748_),
    .C1(_1697_),
    .X(_1749_));
 sky130_fd_sc_hd__mux4_2 _4994_ (.A0(\rf.registers[4][22] ),
    .A1(\rf.registers[5][22] ),
    .A2(\rf.registers[6][22] ),
    .A3(\rf.registers[7][22] ),
    .S0(_1704_),
    .S1(_1707_),
    .X(_1750_));
 sky130_fd_sc_hd__mux4_2 _4995_ (.A0(\rf.registers[0][22] ),
    .A1(\rf.registers[1][22] ),
    .A2(\rf.registers[2][22] ),
    .A3(\rf.registers[3][22] ),
    .S0(_1704_),
    .S1(_1707_),
    .X(_1751_));
 sky130_fd_sc_hd__mux2_2 _4996_ (.A0(_1750_),
    .A1(_1751_),
    .S(_1739_),
    .X(_1752_));
 sky130_fd_sc_hd__a21o_2 _4997_ (.A1(_1717_),
    .A2(_1752_),
    .B1(_1729_),
    .X(_1753_));
 sky130_fd_sc_hd__o22a_2 _4998_ (.A1(_1671_),
    .A2(_1744_),
    .B1(_1749_),
    .B2(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__and2b_2 _4999_ (.A_N(_1639_),
    .B(_1754_),
    .X(_1755_));
 sky130_fd_sc_hd__or2_2 _5000_ (.A(_1668_),
    .B(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__a21bo_2 _5001_ (.A1(_1669_),
    .A2(_1732_),
    .B1_N(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__buf_1 _5002_ (.A(_1639_),
    .X(_1758_));
 sky130_fd_sc_hd__mux4_2 _5003_ (.A0(\rf.registers[20][21] ),
    .A1(\rf.registers[21][21] ),
    .A2(\rf.registers[22][21] ),
    .A3(\rf.registers[23][21] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1759_));
 sky130_fd_sc_hd__mux4_2 _5004_ (.A0(\rf.registers[16][21] ),
    .A1(\rf.registers[17][21] ),
    .A2(\rf.registers[18][21] ),
    .A3(\rf.registers[19][21] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1760_));
 sky130_fd_sc_hd__mux2_2 _5005_ (.A0(_1759_),
    .A1(_1760_),
    .S(_1726_),
    .X(_1761_));
 sky130_fd_sc_hd__mux4_2 _5006_ (.A0(\rf.registers[28][21] ),
    .A1(\rf.registers[29][21] ),
    .A2(\rf.registers[30][21] ),
    .A3(\rf.registers[31][21] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1762_));
 sky130_fd_sc_hd__mux4_2 _5007_ (.A0(\rf.registers[24][21] ),
    .A1(\rf.registers[25][21] ),
    .A2(\rf.registers[26][21] ),
    .A3(\rf.registers[27][21] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1763_));
 sky130_fd_sc_hd__mux2_2 _5008_ (.A0(_1762_),
    .A1(_1763_),
    .S(_1726_),
    .X(_1764_));
 sky130_fd_sc_hd__mux2_2 _5009_ (.A0(_1761_),
    .A1(_1764_),
    .S(_1697_),
    .X(_1765_));
 sky130_fd_sc_hd__buf_1 _5010_ (.A(_1700_),
    .X(_1766_));
 sky130_fd_sc_hd__buf_1 _5011_ (.A(_1704_),
    .X(_1767_));
 sky130_fd_sc_hd__buf_1 _5012_ (.A(_1707_),
    .X(_1768_));
 sky130_fd_sc_hd__mux4_2 _5013_ (.A0(\rf.registers[8][21] ),
    .A1(\rf.registers[9][21] ),
    .A2(\rf.registers[10][21] ),
    .A3(\rf.registers[11][21] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__mux4_2 _5014_ (.A0(\rf.registers[12][21] ),
    .A1(\rf.registers[13][21] ),
    .A2(\rf.registers[14][21] ),
    .A3(\rf.registers[15][21] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1770_));
 sky130_fd_sc_hd__mux2_2 _5015_ (.A0(_1769_),
    .A1(_1770_),
    .S(_1713_),
    .X(_1771_));
 sky130_fd_sc_hd__nand2_2 _5016_ (.A(_1766_),
    .B(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__buf_1 _5017_ (.A(_1717_),
    .X(_1773_));
 sky130_fd_sc_hd__mux4_2 _5018_ (.A0(\rf.registers[4][21] ),
    .A1(\rf.registers[5][21] ),
    .A2(\rf.registers[6][21] ),
    .A3(\rf.registers[7][21] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1774_));
 sky130_fd_sc_hd__mux4_2 _5019_ (.A0(\rf.registers[0][21] ),
    .A1(\rf.registers[1][21] ),
    .A2(\rf.registers[2][21] ),
    .A3(\rf.registers[3][21] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1775_));
 sky130_fd_sc_hd__mux2_2 _5020_ (.A0(_1774_),
    .A1(_1775_),
    .S(_1726_),
    .X(_1776_));
 sky130_fd_sc_hd__buf_1 _5021_ (.A(_1729_),
    .X(_1777_));
 sky130_fd_sc_hd__a21oi_2 _5022_ (.A1(_1773_),
    .A2(_1776_),
    .B1(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__a2bb2o_2 _5023_ (.A1_N(_1672_),
    .A2_N(_1765_),
    .B1(_1772_),
    .B2(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__nor2_2 _5024_ (.A(_1758_),
    .B(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__or2_2 _5025_ (.A(_1168_),
    .B(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__buf_1 _5026_ (.A(_1733_),
    .X(_1782_));
 sky130_fd_sc_hd__mux4_2 _5027_ (.A0(\rf.registers[20][20] ),
    .A1(\rf.registers[21][20] ),
    .A2(\rf.registers[22][20] ),
    .A3(\rf.registers[23][20] ),
    .S0(_1782_),
    .S1(_1680_),
    .X(_1783_));
 sky130_fd_sc_hd__mux4_2 _5028_ (.A0(\rf.registers[16][20] ),
    .A1(\rf.registers[17][20] ),
    .A2(\rf.registers[18][20] ),
    .A3(\rf.registers[19][20] ),
    .S0(_1782_),
    .S1(_1680_),
    .X(_1784_));
 sky130_fd_sc_hd__mux2_2 _5029_ (.A0(_1783_),
    .A1(_1784_),
    .S(_1739_),
    .X(_1785_));
 sky130_fd_sc_hd__mux4_2 _5030_ (.A0(\rf.registers[28][20] ),
    .A1(\rf.registers[29][20] ),
    .A2(\rf.registers[30][20] ),
    .A3(\rf.registers[31][20] ),
    .S0(_1782_),
    .S1(_1680_),
    .X(_1786_));
 sky130_fd_sc_hd__mux4_2 _5031_ (.A0(\rf.registers[24][20] ),
    .A1(\rf.registers[25][20] ),
    .A2(\rf.registers[26][20] ),
    .A3(\rf.registers[27][20] ),
    .S0(_1782_),
    .S1(_1680_),
    .X(_1787_));
 sky130_fd_sc_hd__mux2_2 _5032_ (.A0(_1786_),
    .A1(_1787_),
    .S(_1739_),
    .X(_1788_));
 sky130_fd_sc_hd__mux2_2 _5033_ (.A0(_1785_),
    .A1(_1788_),
    .S(_1699_),
    .X(_1789_));
 sky130_fd_sc_hd__mux4_2 _5034_ (.A0(\rf.registers[8][20] ),
    .A1(\rf.registers[9][20] ),
    .A2(\rf.registers[10][20] ),
    .A3(\rf.registers[11][20] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_1790_));
 sky130_fd_sc_hd__and2_2 _5035_ (.A(_1686_),
    .B(_1790_),
    .X(_1791_));
 sky130_fd_sc_hd__mux4_2 _5036_ (.A0(\rf.registers[12][20] ),
    .A1(\rf.registers[13][20] ),
    .A2(\rf.registers[14][20] ),
    .A3(\rf.registers[15][20] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_1792_));
 sky130_fd_sc_hd__a21o_2 _5037_ (.A1(_1712_),
    .A2(_1792_),
    .B1(_1716_),
    .X(_1793_));
 sky130_fd_sc_hd__mux4_2 _5038_ (.A0(\rf.registers[4][20] ),
    .A1(\rf.registers[5][20] ),
    .A2(\rf.registers[6][20] ),
    .A3(\rf.registers[7][20] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_1794_));
 sky130_fd_sc_hd__mux4_2 _5039_ (.A0(\rf.registers[0][20] ),
    .A1(\rf.registers[1][20] ),
    .A2(\rf.registers[2][20] ),
    .A3(\rf.registers[3][20] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_1795_));
 sky130_fd_sc_hd__mux2_2 _5040_ (.A0(_1794_),
    .A1(_1795_),
    .S(_1739_),
    .X(_1796_));
 sky130_fd_sc_hd__o221a_2 _5041_ (.A1(_1791_),
    .A2(_1793_),
    .B1(_1796_),
    .B2(_1697_),
    .C1(_1671_),
    .X(_1797_));
 sky130_fd_sc_hd__a21oi_2 _5042_ (.A1(_1729_),
    .A2(_1789_),
    .B1(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__buf_1 _5043_ (.A(_1167_),
    .X(_1799_));
 sky130_fd_sc_hd__buf_1 _5044_ (.A(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__o21ai_2 _5045_ (.A1(_1758_),
    .A2(_1798_),
    .B1(_1800_),
    .Y(_1801_));
 sky130_fd_sc_hd__nand2_2 _5046_ (.A(_1781_),
    .B(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__buf_1 _5047_ (.A(_1145_),
    .X(_1803_));
 sky130_fd_sc_hd__mux2_2 _5048_ (.A0(_1757_),
    .A1(_1802_),
    .S(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__mux4_2 _5049_ (.A0(\rf.registers[20][18] ),
    .A1(\rf.registers[21][18] ),
    .A2(\rf.registers[22][18] ),
    .A3(\rf.registers[23][18] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_1805_));
 sky130_fd_sc_hd__mux4_2 _5050_ (.A0(\rf.registers[16][18] ),
    .A1(\rf.registers[17][18] ),
    .A2(\rf.registers[18][18] ),
    .A3(\rf.registers[19][18] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_1806_));
 sky130_fd_sc_hd__mux2_2 _5051_ (.A0(_1805_),
    .A1(_1806_),
    .S(_1739_),
    .X(_1807_));
 sky130_fd_sc_hd__mux4_2 _5052_ (.A0(\rf.registers[28][18] ),
    .A1(\rf.registers[29][18] ),
    .A2(\rf.registers[30][18] ),
    .A3(\rf.registers[31][18] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_1808_));
 sky130_fd_sc_hd__mux4_2 _5053_ (.A0(\rf.registers[24][18] ),
    .A1(\rf.registers[25][18] ),
    .A2(\rf.registers[26][18] ),
    .A3(\rf.registers[27][18] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_1809_));
 sky130_fd_sc_hd__mux2_2 _5054_ (.A0(_1808_),
    .A1(_1809_),
    .S(_1739_),
    .X(_1810_));
 sky130_fd_sc_hd__mux2_2 _5055_ (.A0(_1807_),
    .A1(_1810_),
    .S(_1697_),
    .X(_1811_));
 sky130_fd_sc_hd__mux4_2 _5056_ (.A0(\rf.registers[8][18] ),
    .A1(\rf.registers[9][18] ),
    .A2(\rf.registers[10][18] ),
    .A3(\rf.registers[11][18] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1812_));
 sky130_fd_sc_hd__mux4_2 _5057_ (.A0(\rf.registers[12][18] ),
    .A1(\rf.registers[13][18] ),
    .A2(\rf.registers[14][18] ),
    .A3(\rf.registers[15][18] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1813_));
 sky130_fd_sc_hd__mux2_2 _5058_ (.A0(_1812_),
    .A1(_1813_),
    .S(_1713_),
    .X(_1814_));
 sky130_fd_sc_hd__nand2_2 _5059_ (.A(_1700_),
    .B(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__mux4_2 _5060_ (.A0(\rf.registers[4][18] ),
    .A1(\rf.registers[5][18] ),
    .A2(\rf.registers[6][18] ),
    .A3(\rf.registers[7][18] ),
    .S0(_1704_),
    .S1(_1707_),
    .X(_1816_));
 sky130_fd_sc_hd__mux4_2 _5061_ (.A0(\rf.registers[0][18] ),
    .A1(\rf.registers[1][18] ),
    .A2(\rf.registers[2][18] ),
    .A3(\rf.registers[3][18] ),
    .S0(_1704_),
    .S1(_1707_),
    .X(_1817_));
 sky130_fd_sc_hd__mux2_2 _5062_ (.A0(_1816_),
    .A1(_1817_),
    .S(_1686_),
    .X(_1818_));
 sky130_fd_sc_hd__a21oi_2 _5063_ (.A1(_1717_),
    .A2(_1818_),
    .B1(_1729_),
    .Y(_1819_));
 sky130_fd_sc_hd__a2bb2o_2 _5064_ (.A1_N(_1671_),
    .A2_N(_1811_),
    .B1(_1815_),
    .B2(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__nor2_2 _5065_ (.A(_1758_),
    .B(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__buf_1 _5066_ (.A(_1782_),
    .X(_1822_));
 sky130_fd_sc_hd__buf_1 _5067_ (.A(_1735_),
    .X(_1823_));
 sky130_fd_sc_hd__mux4_2 _5068_ (.A0(\rf.registers[24][19] ),
    .A1(\rf.registers[25][19] ),
    .A2(\rf.registers[26][19] ),
    .A3(\rf.registers[27][19] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__mux4_2 _5069_ (.A0(\rf.registers[28][19] ),
    .A1(\rf.registers[29][19] ),
    .A2(\rf.registers[30][19] ),
    .A3(\rf.registers[31][19] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1825_));
 sky130_fd_sc_hd__mux4_2 _5070_ (.A0(\rf.registers[16][19] ),
    .A1(\rf.registers[17][19] ),
    .A2(\rf.registers[18][19] ),
    .A3(\rf.registers[19][19] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1826_));
 sky130_fd_sc_hd__mux4_2 _5071_ (.A0(\rf.registers[20][19] ),
    .A1(\rf.registers[21][19] ),
    .A2(\rf.registers[22][19] ),
    .A3(\rf.registers[23][19] ),
    .S0(_1676_),
    .S1(_1681_),
    .X(_1827_));
 sky130_fd_sc_hd__buf_1 _5072_ (.A(_1716_),
    .X(_1828_));
 sky130_fd_sc_hd__mux4_2 _5073_ (.A0(_1824_),
    .A1(_1825_),
    .A2(_1826_),
    .A3(_1827_),
    .S0(_1713_),
    .S1(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__mux4_2 _5074_ (.A0(\rf.registers[12][19] ),
    .A1(\rf.registers[13][19] ),
    .A2(\rf.registers[14][19] ),
    .A3(\rf.registers[15][19] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1830_));
 sky130_fd_sc_hd__mux4_2 _5075_ (.A0(\rf.registers[8][19] ),
    .A1(\rf.registers[9][19] ),
    .A2(\rf.registers[10][19] ),
    .A3(\rf.registers[11][19] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1831_));
 sky130_fd_sc_hd__mux2_2 _5076_ (.A0(_1830_),
    .A1(_1831_),
    .S(_1686_),
    .X(_1832_));
 sky130_fd_sc_hd__nand2_2 _5077_ (.A(_1700_),
    .B(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__mux4_2 _5078_ (.A0(\rf.registers[4][19] ),
    .A1(\rf.registers[5][19] ),
    .A2(\rf.registers[6][19] ),
    .A3(\rf.registers[7][19] ),
    .S0(_1704_),
    .S1(_1707_),
    .X(_1834_));
 sky130_fd_sc_hd__mux4_2 _5079_ (.A0(\rf.registers[0][19] ),
    .A1(\rf.registers[1][19] ),
    .A2(\rf.registers[2][19] ),
    .A3(\rf.registers[3][19] ),
    .S0(_1704_),
    .S1(_1707_),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_2 _5080_ (.A0(_1834_),
    .A1(_1835_),
    .S(_1686_),
    .X(_1836_));
 sky130_fd_sc_hd__a21oi_2 _5081_ (.A1(_1717_),
    .A2(_1836_),
    .B1(_1729_),
    .Y(_1837_));
 sky130_fd_sc_hd__a2bb2o_2 _5082_ (.A1_N(_1671_),
    .A2_N(_1829_),
    .B1(_1833_),
    .B2(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__buf_1 _5083_ (.A(_1667_),
    .X(_1839_));
 sky130_fd_sc_hd__o21a_2 _5084_ (.A1(_1758_),
    .A2(_1838_),
    .B1(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__o21bai_2 _5085_ (.A1(_1669_),
    .A2(_1821_),
    .B1_N(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__buf_1 _5086_ (.A(_1638_),
    .X(_1842_));
 sky130_fd_sc_hd__mux4_2 _5087_ (.A0(\rf.registers[20][17] ),
    .A1(\rf.registers[21][17] ),
    .A2(\rf.registers[22][17] ),
    .A3(\rf.registers[23][17] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1843_));
 sky130_fd_sc_hd__mux4_2 _5088_ (.A0(\rf.registers[16][17] ),
    .A1(\rf.registers[17][17] ),
    .A2(\rf.registers[18][17] ),
    .A3(\rf.registers[19][17] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1844_));
 sky130_fd_sc_hd__mux2_2 _5089_ (.A0(_1843_),
    .A1(_1844_),
    .S(_1686_),
    .X(_1845_));
 sky130_fd_sc_hd__mux4_2 _5090_ (.A0(\rf.registers[28][17] ),
    .A1(\rf.registers[29][17] ),
    .A2(\rf.registers[30][17] ),
    .A3(\rf.registers[31][17] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1846_));
 sky130_fd_sc_hd__mux4_2 _5091_ (.A0(\rf.registers[24][17] ),
    .A1(\rf.registers[25][17] ),
    .A2(\rf.registers[26][17] ),
    .A3(\rf.registers[27][17] ),
    .S0(_1689_),
    .S1(_1693_),
    .X(_1847_));
 sky130_fd_sc_hd__mux2_2 _5092_ (.A0(_1846_),
    .A1(_1847_),
    .S(_1686_),
    .X(_1848_));
 sky130_fd_sc_hd__mux2_2 _5093_ (.A0(_1845_),
    .A1(_1848_),
    .S(_1697_),
    .X(_1849_));
 sky130_fd_sc_hd__mux4_2 _5094_ (.A0(\rf.registers[8][17] ),
    .A1(\rf.registers[9][17] ),
    .A2(\rf.registers[10][17] ),
    .A3(\rf.registers[11][17] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1850_));
 sky130_fd_sc_hd__mux4_2 _5095_ (.A0(\rf.registers[12][17] ),
    .A1(\rf.registers[13][17] ),
    .A2(\rf.registers[14][17] ),
    .A3(\rf.registers[15][17] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1851_));
 sky130_fd_sc_hd__mux2_2 _5096_ (.A0(_1850_),
    .A1(_1851_),
    .S(_1713_),
    .X(_1852_));
 sky130_fd_sc_hd__nand2_2 _5097_ (.A(_1700_),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__mux4_2 _5098_ (.A0(\rf.registers[4][17] ),
    .A1(\rf.registers[5][17] ),
    .A2(\rf.registers[6][17] ),
    .A3(\rf.registers[7][17] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_1854_));
 sky130_fd_sc_hd__mux4_2 _5099_ (.A0(\rf.registers[0][17] ),
    .A1(\rf.registers[1][17] ),
    .A2(\rf.registers[2][17] ),
    .A3(\rf.registers[3][17] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_1855_));
 sky130_fd_sc_hd__mux2_2 _5100_ (.A0(_1854_),
    .A1(_1855_),
    .S(_1726_),
    .X(_1856_));
 sky130_fd_sc_hd__a21oi_2 _5101_ (.A1(_1717_),
    .A2(_1856_),
    .B1(_1729_),
    .Y(_1857_));
 sky130_fd_sc_hd__a2bb2o_2 _5102_ (.A1_N(_1672_),
    .A2_N(_1849_),
    .B1(_1853_),
    .B2(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__nor2_2 _5103_ (.A(_1842_),
    .B(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__or2_2 _5104_ (.A(_1168_),
    .B(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__mux4_2 _5105_ (.A0(\rf.registers[24][16] ),
    .A1(\rf.registers[25][16] ),
    .A2(\rf.registers[26][16] ),
    .A3(\rf.registers[27][16] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1861_));
 sky130_fd_sc_hd__mux4_2 _5106_ (.A0(\rf.registers[28][16] ),
    .A1(\rf.registers[29][16] ),
    .A2(\rf.registers[30][16] ),
    .A3(\rf.registers[31][16] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1862_));
 sky130_fd_sc_hd__mux4_2 _5107_ (.A0(\rf.registers[16][16] ),
    .A1(\rf.registers[17][16] ),
    .A2(\rf.registers[18][16] ),
    .A3(\rf.registers[19][16] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1863_));
 sky130_fd_sc_hd__mux4_2 _5108_ (.A0(\rf.registers[20][16] ),
    .A1(\rf.registers[21][16] ),
    .A2(\rf.registers[22][16] ),
    .A3(\rf.registers[23][16] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1864_));
 sky130_fd_sc_hd__mux4_2 _5109_ (.A0(_1861_),
    .A1(_1862_),
    .A2(_1863_),
    .A3(_1864_),
    .S0(_1713_),
    .S1(_1717_),
    .X(_1865_));
 sky130_fd_sc_hd__mux4_2 _5110_ (.A0(\rf.registers[8][16] ),
    .A1(\rf.registers[9][16] ),
    .A2(\rf.registers[10][16] ),
    .A3(\rf.registers[11][16] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1866_));
 sky130_fd_sc_hd__mux4_2 _5111_ (.A0(\rf.registers[12][16] ),
    .A1(\rf.registers[13][16] ),
    .A2(\rf.registers[14][16] ),
    .A3(\rf.registers[15][16] ),
    .S0(_1720_),
    .S1(_1723_),
    .X(_1867_));
 sky130_fd_sc_hd__mux2_2 _5112_ (.A0(_1866_),
    .A1(_1867_),
    .S(_1713_),
    .X(_1868_));
 sky130_fd_sc_hd__nor2_2 _5113_ (.A(_1717_),
    .B(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__mux4_2 _5114_ (.A0(\rf.registers[4][16] ),
    .A1(\rf.registers[5][16] ),
    .A2(\rf.registers[6][16] ),
    .A3(\rf.registers[7][16] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_1870_));
 sky130_fd_sc_hd__mux4_2 _5115_ (.A0(\rf.registers[0][16] ),
    .A1(\rf.registers[1][16] ),
    .A2(\rf.registers[2][16] ),
    .A3(\rf.registers[3][16] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_1871_));
 sky130_fd_sc_hd__mux2_2 _5116_ (.A0(_1870_),
    .A1(_1871_),
    .S(_1726_),
    .X(_1872_));
 sky130_fd_sc_hd__o21ai_2 _5117_ (.A1(_1700_),
    .A2(_1872_),
    .B1(_1671_),
    .Y(_1873_));
 sky130_fd_sc_hd__o2bb2a_2 _5118_ (.A1_N(_1777_),
    .A2_N(_1865_),
    .B1(_1869_),
    .B2(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__o21ai_2 _5119_ (.A1(_1758_),
    .A2(_1874_),
    .B1(_1800_),
    .Y(_1875_));
 sky130_fd_sc_hd__nand2_2 _5120_ (.A(_1860_),
    .B(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__buf_1 _5121_ (.A(_1145_),
    .X(_1877_));
 sky130_fd_sc_hd__mux2_2 _5122_ (.A0(_1841_),
    .A1(_1876_),
    .S(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__buf_1 _5123_ (.A(_1126_),
    .X(_1879_));
 sky130_fd_sc_hd__mux2_2 _5124_ (.A0(_1804_),
    .A1(_1878_),
    .S(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__buf_1 _5125_ (.A(_1720_),
    .X(_1881_));
 sky130_fd_sc_hd__buf_1 _5126_ (.A(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__buf_1 _5127_ (.A(_1723_),
    .X(_1883_));
 sky130_fd_sc_hd__buf_1 _5128_ (.A(_1883_),
    .X(_1884_));
 sky130_fd_sc_hd__mux4_2 _5129_ (.A0(\rf.registers[24][31] ),
    .A1(\rf.registers[25][31] ),
    .A2(\rf.registers[26][31] ),
    .A3(\rf.registers[27][31] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__mux4_2 _5130_ (.A0(\rf.registers[28][31] ),
    .A1(\rf.registers[29][31] ),
    .A2(\rf.registers[30][31] ),
    .A3(\rf.registers[31][31] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1886_));
 sky130_fd_sc_hd__mux4_2 _5131_ (.A0(\rf.registers[16][31] ),
    .A1(\rf.registers[17][31] ),
    .A2(\rf.registers[18][31] ),
    .A3(\rf.registers[19][31] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1887_));
 sky130_fd_sc_hd__mux4_2 _5132_ (.A0(\rf.registers[20][31] ),
    .A1(\rf.registers[21][31] ),
    .A2(\rf.registers[22][31] ),
    .A3(\rf.registers[23][31] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1888_));
 sky130_fd_sc_hd__buf_1 _5133_ (.A(_1713_),
    .X(_1889_));
 sky130_fd_sc_hd__mux4_2 _5134_ (.A0(_1885_),
    .A1(_1886_),
    .A2(_1887_),
    .A3(_1888_),
    .S0(_1889_),
    .S1(_1773_),
    .X(_1890_));
 sky130_fd_sc_hd__mux4_2 _5135_ (.A0(\rf.registers[8][31] ),
    .A1(\rf.registers[9][31] ),
    .A2(\rf.registers[10][31] ),
    .A3(\rf.registers[11][31] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1891_));
 sky130_fd_sc_hd__mux4_2 _5136_ (.A0(\rf.registers[12][31] ),
    .A1(\rf.registers[13][31] ),
    .A2(\rf.registers[14][31] ),
    .A3(\rf.registers[15][31] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1892_));
 sky130_fd_sc_hd__mux2_2 _5137_ (.A0(_1891_),
    .A1(_1892_),
    .S(_1889_),
    .X(_1893_));
 sky130_fd_sc_hd__nor2_2 _5138_ (.A(_1773_),
    .B(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__buf_1 _5139_ (.A(_1689_),
    .X(_1895_));
 sky130_fd_sc_hd__buf_1 _5140_ (.A(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__buf_1 _5141_ (.A(_1693_),
    .X(_1897_));
 sky130_fd_sc_hd__buf_1 _5142_ (.A(_1897_),
    .X(_1898_));
 sky130_fd_sc_hd__mux4_2 _5143_ (.A0(\rf.registers[4][31] ),
    .A1(\rf.registers[5][31] ),
    .A2(\rf.registers[6][31] ),
    .A3(\rf.registers[7][31] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__mux4_2 _5144_ (.A0(\rf.registers[0][31] ),
    .A1(\rf.registers[1][31] ),
    .A2(\rf.registers[2][31] ),
    .A3(\rf.registers[3][31] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1900_));
 sky130_fd_sc_hd__buf_1 _5145_ (.A(_1726_),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_2 _5146_ (.A0(_1899_),
    .A1(_1900_),
    .S(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__o21ai_2 _5147_ (.A1(_1766_),
    .A2(_1902_),
    .B1(_1672_),
    .Y(_1903_));
 sky130_fd_sc_hd__o2bb2a_2 _5148_ (.A1_N(_1777_),
    .A2_N(_1890_),
    .B1(_1894_),
    .B2(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__nor2_2 _5149_ (.A(_1842_),
    .B(_1904_),
    .Y(_1905_));
 sky130_fd_sc_hd__mux4_2 _5150_ (.A0(\rf.registers[20][30] ),
    .A1(\rf.registers[21][30] ),
    .A2(\rf.registers[22][30] ),
    .A3(\rf.registers[23][30] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_1906_));
 sky130_fd_sc_hd__mux4_2 _5151_ (.A0(\rf.registers[16][30] ),
    .A1(\rf.registers[17][30] ),
    .A2(\rf.registers[18][30] ),
    .A3(\rf.registers[19][30] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_1907_));
 sky130_fd_sc_hd__mux2_2 _5152_ (.A0(_1906_),
    .A1(_1907_),
    .S(_1745_),
    .X(_1908_));
 sky130_fd_sc_hd__mux4_2 _5153_ (.A0(\rf.registers[28][30] ),
    .A1(\rf.registers[29][30] ),
    .A2(\rf.registers[30][30] ),
    .A3(\rf.registers[31][30] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_1909_));
 sky130_fd_sc_hd__mux4_2 _5154_ (.A0(\rf.registers[24][30] ),
    .A1(\rf.registers[25][30] ),
    .A2(\rf.registers[26][30] ),
    .A3(\rf.registers[27][30] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_1910_));
 sky130_fd_sc_hd__mux2_2 _5155_ (.A0(_1909_),
    .A1(_1910_),
    .S(_1745_),
    .X(_1911_));
 sky130_fd_sc_hd__mux2_2 _5156_ (.A0(_1908_),
    .A1(_1911_),
    .S(_1700_),
    .X(_1912_));
 sky130_fd_sc_hd__mux4_2 _5157_ (.A0(\rf.registers[8][30] ),
    .A1(\rf.registers[9][30] ),
    .A2(\rf.registers[10][30] ),
    .A3(\rf.registers[11][30] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_1913_));
 sky130_fd_sc_hd__mux4_2 _5158_ (.A0(\rf.registers[12][30] ),
    .A1(\rf.registers[13][30] ),
    .A2(\rf.registers[14][30] ),
    .A3(\rf.registers[15][30] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_2 _5159_ (.A0(_1913_),
    .A1(_1914_),
    .S(_1889_),
    .X(_1915_));
 sky130_fd_sc_hd__nor2_2 _5160_ (.A(_1773_),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__mux4_2 _5161_ (.A0(\rf.registers[4][30] ),
    .A1(\rf.registers[5][30] ),
    .A2(\rf.registers[6][30] ),
    .A3(\rf.registers[7][30] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_1917_));
 sky130_fd_sc_hd__buf_1 _5162_ (.A(_1822_),
    .X(_1918_));
 sky130_fd_sc_hd__buf_1 _5163_ (.A(_1823_),
    .X(_1919_));
 sky130_fd_sc_hd__mux4_2 _5164_ (.A0(\rf.registers[0][30] ),
    .A1(\rf.registers[1][30] ),
    .A2(\rf.registers[2][30] ),
    .A3(\rf.registers[3][30] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__mux2_2 _5165_ (.A0(_1917_),
    .A1(_1920_),
    .S(_1901_),
    .X(_1921_));
 sky130_fd_sc_hd__o21ai_2 _5166_ (.A1(_1766_),
    .A2(_1921_),
    .B1(_1672_),
    .Y(_1922_));
 sky130_fd_sc_hd__o2bb2a_2 _5167_ (.A1_N(_1777_),
    .A2_N(_1912_),
    .B1(_1916_),
    .B2(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__or2_2 _5168_ (.A(_1639_),
    .B(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__nand2_2 _5169_ (.A(_1169_),
    .B(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__o21ai_2 _5170_ (.A1(_1169_),
    .A2(_1905_),
    .B1(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__mux4_2 _5171_ (.A0(\rf.registers[20][29] ),
    .A1(\rf.registers[21][29] ),
    .A2(\rf.registers[22][29] ),
    .A3(\rf.registers[23][29] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1927_));
 sky130_fd_sc_hd__mux4_2 _5172_ (.A0(\rf.registers[16][29] ),
    .A1(\rf.registers[17][29] ),
    .A2(\rf.registers[18][29] ),
    .A3(\rf.registers[19][29] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1928_));
 sky130_fd_sc_hd__mux2_2 _5173_ (.A0(_1927_),
    .A1(_1928_),
    .S(_1745_),
    .X(_1929_));
 sky130_fd_sc_hd__mux4_2 _5174_ (.A0(\rf.registers[28][29] ),
    .A1(\rf.registers[29][29] ),
    .A2(\rf.registers[30][29] ),
    .A3(\rf.registers[31][29] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1930_));
 sky130_fd_sc_hd__mux4_2 _5175_ (.A0(\rf.registers[24][29] ),
    .A1(\rf.registers[25][29] ),
    .A2(\rf.registers[26][29] ),
    .A3(\rf.registers[27][29] ),
    .S0(_1705_),
    .S1(_1708_),
    .X(_1931_));
 sky130_fd_sc_hd__mux2_2 _5176_ (.A0(_1930_),
    .A1(_1931_),
    .S(_1726_),
    .X(_1932_));
 sky130_fd_sc_hd__mux2_2 _5177_ (.A0(_1929_),
    .A1(_1932_),
    .S(_1700_),
    .X(_1933_));
 sky130_fd_sc_hd__mux4_2 _5178_ (.A0(\rf.registers[4][29] ),
    .A1(\rf.registers[5][29] ),
    .A2(\rf.registers[6][29] ),
    .A3(\rf.registers[7][29] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1934_));
 sky130_fd_sc_hd__and2_2 _5179_ (.A(_1889_),
    .B(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__mux4_2 _5180_ (.A0(\rf.registers[0][29] ),
    .A1(\rf.registers[1][29] ),
    .A2(\rf.registers[2][29] ),
    .A3(\rf.registers[3][29] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_1936_));
 sky130_fd_sc_hd__a21o_2 _5181_ (.A1(_1745_),
    .A2(_1936_),
    .B1(_1697_),
    .X(_1937_));
 sky130_fd_sc_hd__mux4_2 _5182_ (.A0(\rf.registers[8][29] ),
    .A1(\rf.registers[9][29] ),
    .A2(\rf.registers[10][29] ),
    .A3(\rf.registers[11][29] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1938_));
 sky130_fd_sc_hd__mux4_2 _5183_ (.A0(\rf.registers[12][29] ),
    .A1(\rf.registers[13][29] ),
    .A2(\rf.registers[14][29] ),
    .A3(\rf.registers[15][29] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_2 _5184_ (.A0(_1938_),
    .A1(_1939_),
    .S(_1713_),
    .X(_1940_));
 sky130_fd_sc_hd__o221a_2 _5185_ (.A1(_1935_),
    .A2(_1937_),
    .B1(_1940_),
    .B2(_1773_),
    .C1(_1671_),
    .X(_1941_));
 sky130_fd_sc_hd__a21o_2 _5186_ (.A1(_1777_),
    .A2(_1933_),
    .B1(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__and2b_2 _5187_ (.A_N(_1638_),
    .B(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__nor2_2 _5188_ (.A(_1800_),
    .B(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__mux4_2 _5189_ (.A0(\rf.registers[24][28] ),
    .A1(\rf.registers[25][28] ),
    .A2(\rf.registers[26][28] ),
    .A3(\rf.registers[27][28] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1945_));
 sky130_fd_sc_hd__mux4_2 _5190_ (.A0(\rf.registers[28][28] ),
    .A1(\rf.registers[29][28] ),
    .A2(\rf.registers[30][28] ),
    .A3(\rf.registers[31][28] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1946_));
 sky130_fd_sc_hd__mux4_2 _5191_ (.A0(\rf.registers[16][28] ),
    .A1(\rf.registers[17][28] ),
    .A2(\rf.registers[18][28] ),
    .A3(\rf.registers[19][28] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1947_));
 sky130_fd_sc_hd__mux4_2 _5192_ (.A0(\rf.registers[20][28] ),
    .A1(\rf.registers[21][28] ),
    .A2(\rf.registers[22][28] ),
    .A3(\rf.registers[23][28] ),
    .S0(_1882_),
    .S1(_1884_),
    .X(_1948_));
 sky130_fd_sc_hd__mux4_2 _5193_ (.A0(_1945_),
    .A1(_1946_),
    .A2(_1947_),
    .A3(_1948_),
    .S0(_1889_),
    .S1(_1773_),
    .X(_1949_));
 sky130_fd_sc_hd__mux4_2 _5194_ (.A0(\rf.registers[4][28] ),
    .A1(\rf.registers[5][28] ),
    .A2(\rf.registers[6][28] ),
    .A3(\rf.registers[7][28] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1950_));
 sky130_fd_sc_hd__and2_2 _5195_ (.A(_1889_),
    .B(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__mux4_2 _5196_ (.A0(\rf.registers[0][28] ),
    .A1(\rf.registers[1][28] ),
    .A2(\rf.registers[2][28] ),
    .A3(\rf.registers[3][28] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1952_));
 sky130_fd_sc_hd__a21o_2 _5197_ (.A1(_1901_),
    .A2(_1952_),
    .B1(_1766_),
    .X(_1953_));
 sky130_fd_sc_hd__mux4_2 _5198_ (.A0(\rf.registers[8][28] ),
    .A1(\rf.registers[9][28] ),
    .A2(\rf.registers[10][28] ),
    .A3(\rf.registers[11][28] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1954_));
 sky130_fd_sc_hd__mux4_2 _5199_ (.A0(\rf.registers[12][28] ),
    .A1(\rf.registers[13][28] ),
    .A2(\rf.registers[14][28] ),
    .A3(\rf.registers[15][28] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1955_));
 sky130_fd_sc_hd__mux2_2 _5200_ (.A0(_1954_),
    .A1(_1955_),
    .S(_1889_),
    .X(_1956_));
 sky130_fd_sc_hd__o221a_2 _5201_ (.A1(_1951_),
    .A2(_1953_),
    .B1(_1956_),
    .B2(_1773_),
    .C1(_1672_),
    .X(_1957_));
 sky130_fd_sc_hd__a21oi_2 _5202_ (.A1(_1777_),
    .A2(_1949_),
    .B1(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__nor2_2 _5203_ (.A(_1842_),
    .B(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__nor2_2 _5204_ (.A(_1839_),
    .B(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hd__or2_2 _5205_ (.A(_1944_),
    .B(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__mux2_2 _5206_ (.A0(_1926_),
    .A1(_1961_),
    .S(_1877_),
    .X(_1962_));
 sky130_fd_sc_hd__mux4_2 _5207_ (.A0(\rf.registers[20][27] ),
    .A1(\rf.registers[21][27] ),
    .A2(\rf.registers[22][27] ),
    .A3(\rf.registers[23][27] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1963_));
 sky130_fd_sc_hd__mux4_2 _5208_ (.A0(\rf.registers[16][27] ),
    .A1(\rf.registers[17][27] ),
    .A2(\rf.registers[18][27] ),
    .A3(\rf.registers[19][27] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1964_));
 sky130_fd_sc_hd__mux2_2 _5209_ (.A0(_1963_),
    .A1(_1964_),
    .S(_1745_),
    .X(_1965_));
 sky130_fd_sc_hd__mux4_2 _5210_ (.A0(\rf.registers[28][27] ),
    .A1(\rf.registers[29][27] ),
    .A2(\rf.registers[30][27] ),
    .A3(\rf.registers[31][27] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1966_));
 sky130_fd_sc_hd__mux4_2 _5211_ (.A0(\rf.registers[24][27] ),
    .A1(\rf.registers[25][27] ),
    .A2(\rf.registers[26][27] ),
    .A3(\rf.registers[27][27] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_1967_));
 sky130_fd_sc_hd__mux2_2 _5212_ (.A0(_1966_),
    .A1(_1967_),
    .S(_1745_),
    .X(_1968_));
 sky130_fd_sc_hd__mux2_2 _5213_ (.A0(_1965_),
    .A1(_1968_),
    .S(_1700_),
    .X(_1969_));
 sky130_fd_sc_hd__mux4_2 _5214_ (.A0(\rf.registers[8][27] ),
    .A1(\rf.registers[9][27] ),
    .A2(\rf.registers[10][27] ),
    .A3(\rf.registers[11][27] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_1970_));
 sky130_fd_sc_hd__mux4_2 _5215_ (.A0(\rf.registers[12][27] ),
    .A1(\rf.registers[13][27] ),
    .A2(\rf.registers[14][27] ),
    .A3(\rf.registers[15][27] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_1971_));
 sky130_fd_sc_hd__mux2_2 _5216_ (.A0(_1970_),
    .A1(_1971_),
    .S(_1889_),
    .X(_1972_));
 sky130_fd_sc_hd__nor2_2 _5217_ (.A(_1773_),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__mux4_2 _5218_ (.A0(\rf.registers[4][27] ),
    .A1(\rf.registers[5][27] ),
    .A2(\rf.registers[6][27] ),
    .A3(\rf.registers[7][27] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_1974_));
 sky130_fd_sc_hd__mux4_2 _5219_ (.A0(\rf.registers[0][27] ),
    .A1(\rf.registers[1][27] ),
    .A2(\rf.registers[2][27] ),
    .A3(\rf.registers[3][27] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_1975_));
 sky130_fd_sc_hd__mux2_2 _5220_ (.A0(_1974_),
    .A1(_1975_),
    .S(_1745_),
    .X(_1976_));
 sky130_fd_sc_hd__o21ai_2 _5221_ (.A1(_1766_),
    .A2(_1976_),
    .B1(_1672_),
    .Y(_1977_));
 sky130_fd_sc_hd__o2bb2a_2 _5222_ (.A1_N(_1777_),
    .A2_N(_1969_),
    .B1(_1973_),
    .B2(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__nor2_2 _5223_ (.A(_1842_),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__nor2_2 _5224_ (.A(_1800_),
    .B(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__mux4_2 _5225_ (.A0(\rf.registers[20][26] ),
    .A1(\rf.registers[21][26] ),
    .A2(\rf.registers[22][26] ),
    .A3(\rf.registers[23][26] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_1981_));
 sky130_fd_sc_hd__mux4_2 _5226_ (.A0(\rf.registers[16][26] ),
    .A1(\rf.registers[17][26] ),
    .A2(\rf.registers[18][26] ),
    .A3(\rf.registers[19][26] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_1982_));
 sky130_fd_sc_hd__mux2_2 _5227_ (.A0(_1981_),
    .A1(_1982_),
    .S(_1901_),
    .X(_1983_));
 sky130_fd_sc_hd__mux4_2 _5228_ (.A0(\rf.registers[28][26] ),
    .A1(\rf.registers[29][26] ),
    .A2(\rf.registers[30][26] ),
    .A3(\rf.registers[31][26] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_1984_));
 sky130_fd_sc_hd__mux4_2 _5229_ (.A0(\rf.registers[24][26] ),
    .A1(\rf.registers[25][26] ),
    .A2(\rf.registers[26][26] ),
    .A3(\rf.registers[27][26] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_1985_));
 sky130_fd_sc_hd__mux2_2 _5230_ (.A0(_1984_),
    .A1(_1985_),
    .S(_1901_),
    .X(_1986_));
 sky130_fd_sc_hd__mux2_2 _5231_ (.A0(_1983_),
    .A1(_1986_),
    .S(_1766_),
    .X(_1987_));
 sky130_fd_sc_hd__mux4_2 _5232_ (.A0(\rf.registers[12][26] ),
    .A1(\rf.registers[13][26] ),
    .A2(\rf.registers[14][26] ),
    .A3(\rf.registers[15][26] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1988_));
 sky130_fd_sc_hd__mux4_2 _5233_ (.A0(\rf.registers[8][26] ),
    .A1(\rf.registers[9][26] ),
    .A2(\rf.registers[10][26] ),
    .A3(\rf.registers[11][26] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1989_));
 sky130_fd_sc_hd__mux2_2 _5234_ (.A0(_1988_),
    .A1(_1989_),
    .S(_1901_),
    .X(_1990_));
 sky130_fd_sc_hd__mux4_2 _5235_ (.A0(\rf.registers[4][26] ),
    .A1(\rf.registers[5][26] ),
    .A2(\rf.registers[6][26] ),
    .A3(\rf.registers[7][26] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1991_));
 sky130_fd_sc_hd__and2_2 _5236_ (.A(_1889_),
    .B(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__mux4_2 _5237_ (.A0(\rf.registers[0][26] ),
    .A1(\rf.registers[1][26] ),
    .A2(\rf.registers[2][26] ),
    .A3(\rf.registers[3][26] ),
    .S0(_1896_),
    .S1(_1898_),
    .X(_1993_));
 sky130_fd_sc_hd__a21o_2 _5238_ (.A1(_1901_),
    .A2(_1993_),
    .B1(_1766_),
    .X(_1994_));
 sky130_fd_sc_hd__o221a_2 _5239_ (.A1(_1773_),
    .A2(_1990_),
    .B1(_1992_),
    .B2(_1994_),
    .C1(_1672_),
    .X(_1995_));
 sky130_fd_sc_hd__a21oi_2 _5240_ (.A1(_1777_),
    .A2(_1987_),
    .B1(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__nor2_2 _5241_ (.A(_1842_),
    .B(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__nor2_2 _5242_ (.A(_1839_),
    .B(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__or2_2 _5243_ (.A(_1980_),
    .B(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__mux4_2 _5244_ (.A0(\rf.registers[20][25] ),
    .A1(\rf.registers[21][25] ),
    .A2(\rf.registers[22][25] ),
    .A3(\rf.registers[23][25] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_2000_));
 sky130_fd_sc_hd__mux4_2 _5245_ (.A0(\rf.registers[16][25] ),
    .A1(\rf.registers[17][25] ),
    .A2(\rf.registers[18][25] ),
    .A3(\rf.registers[19][25] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_2001_));
 sky130_fd_sc_hd__mux2_2 _5246_ (.A0(_2000_),
    .A1(_2001_),
    .S(_1726_),
    .X(_2002_));
 sky130_fd_sc_hd__mux4_2 _5247_ (.A0(\rf.registers[28][25] ),
    .A1(\rf.registers[29][25] ),
    .A2(\rf.registers[30][25] ),
    .A3(\rf.registers[31][25] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_2003_));
 sky130_fd_sc_hd__mux4_2 _5248_ (.A0(\rf.registers[24][25] ),
    .A1(\rf.registers[25][25] ),
    .A2(\rf.registers[26][25] ),
    .A3(\rf.registers[27][25] ),
    .S0(_1822_),
    .S1(_1823_),
    .X(_2004_));
 sky130_fd_sc_hd__mux2_2 _5249_ (.A0(_2003_),
    .A1(_2004_),
    .S(_1726_),
    .X(_2005_));
 sky130_fd_sc_hd__mux2_2 _5250_ (.A0(_2002_),
    .A1(_2005_),
    .S(_1700_),
    .X(_2006_));
 sky130_fd_sc_hd__mux4_2 _5251_ (.A0(\rf.registers[8][25] ),
    .A1(\rf.registers[9][25] ),
    .A2(\rf.registers[10][25] ),
    .A3(\rf.registers[11][25] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_2007_));
 sky130_fd_sc_hd__mux4_2 _5252_ (.A0(\rf.registers[12][25] ),
    .A1(\rf.registers[13][25] ),
    .A2(\rf.registers[14][25] ),
    .A3(\rf.registers[15][25] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_2008_));
 sky130_fd_sc_hd__mux2_2 _5253_ (.A0(_2007_),
    .A1(_2008_),
    .S(_1713_),
    .X(_2009_));
 sky130_fd_sc_hd__nor2_2 _5254_ (.A(_1773_),
    .B(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__mux4_2 _5255_ (.A0(\rf.registers[4][25] ),
    .A1(\rf.registers[5][25] ),
    .A2(\rf.registers[6][25] ),
    .A3(\rf.registers[7][25] ),
    .S0(_1895_),
    .S1(_1897_),
    .X(_2011_));
 sky130_fd_sc_hd__mux4_2 _5256_ (.A0(\rf.registers[0][25] ),
    .A1(\rf.registers[1][25] ),
    .A2(\rf.registers[2][25] ),
    .A3(\rf.registers[3][25] ),
    .S0(_1767_),
    .S1(_1768_),
    .X(_2012_));
 sky130_fd_sc_hd__mux2_2 _5257_ (.A0(_2011_),
    .A1(_2012_),
    .S(_1745_),
    .X(_2013_));
 sky130_fd_sc_hd__o21ai_2 _5258_ (.A1(_1766_),
    .A2(_2013_),
    .B1(_1672_),
    .Y(_2014_));
 sky130_fd_sc_hd__o2bb2a_2 _5259_ (.A1_N(_1777_),
    .A2_N(_2006_),
    .B1(_2010_),
    .B2(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__or2_2 _5260_ (.A(_1638_),
    .B(_2015_),
    .X(_2016_));
 sky130_fd_sc_hd__and2_2 _5261_ (.A(_1668_),
    .B(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__mux4_2 _5262_ (.A0(\rf.registers[20][24] ),
    .A1(\rf.registers[21][24] ),
    .A2(\rf.registers[22][24] ),
    .A3(\rf.registers[23][24] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_2018_));
 sky130_fd_sc_hd__mux4_2 _5263_ (.A0(\rf.registers[16][24] ),
    .A1(\rf.registers[17][24] ),
    .A2(\rf.registers[18][24] ),
    .A3(\rf.registers[19][24] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_2019_));
 sky130_fd_sc_hd__mux2_2 _5264_ (.A0(_2018_),
    .A1(_2019_),
    .S(_1901_),
    .X(_2020_));
 sky130_fd_sc_hd__mux4_2 _5265_ (.A0(\rf.registers[28][24] ),
    .A1(\rf.registers[29][24] ),
    .A2(\rf.registers[30][24] ),
    .A3(\rf.registers[31][24] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_2021_));
 sky130_fd_sc_hd__mux4_2 _5266_ (.A0(\rf.registers[24][24] ),
    .A1(\rf.registers[25][24] ),
    .A2(\rf.registers[26][24] ),
    .A3(\rf.registers[27][24] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_2022_));
 sky130_fd_sc_hd__mux2_2 _5267_ (.A0(_2021_),
    .A1(_2022_),
    .S(_1745_),
    .X(_2023_));
 sky130_fd_sc_hd__mux2_2 _5268_ (.A0(_2020_),
    .A1(_2023_),
    .S(_1766_),
    .X(_2024_));
 sky130_fd_sc_hd__mux4_2 _5269_ (.A0(\rf.registers[12][24] ),
    .A1(\rf.registers[13][24] ),
    .A2(\rf.registers[14][24] ),
    .A3(\rf.registers[15][24] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_2025_));
 sky130_fd_sc_hd__and2_2 _5270_ (.A(_1889_),
    .B(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__mux4_2 _5271_ (.A0(\rf.registers[8][24] ),
    .A1(\rf.registers[9][24] ),
    .A2(\rf.registers[10][24] ),
    .A3(\rf.registers[11][24] ),
    .S0(_1881_),
    .S1(_1883_),
    .X(_2027_));
 sky130_fd_sc_hd__a21o_2 _5272_ (.A1(_1901_),
    .A2(_2027_),
    .B1(_1717_),
    .X(_2028_));
 sky130_fd_sc_hd__mux4_2 _5273_ (.A0(\rf.registers[4][24] ),
    .A1(\rf.registers[5][24] ),
    .A2(\rf.registers[6][24] ),
    .A3(\rf.registers[7][24] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_2029_));
 sky130_fd_sc_hd__mux4_2 _5274_ (.A0(\rf.registers[0][24] ),
    .A1(\rf.registers[1][24] ),
    .A2(\rf.registers[2][24] ),
    .A3(\rf.registers[3][24] ),
    .S0(_1918_),
    .S1(_1919_),
    .X(_2030_));
 sky130_fd_sc_hd__mux2_2 _5275_ (.A0(_2029_),
    .A1(_2030_),
    .S(_1901_),
    .X(_2031_));
 sky130_fd_sc_hd__o221a_2 _5276_ (.A1(_2026_),
    .A2(_2028_),
    .B1(_2031_),
    .B2(_1766_),
    .C1(_1672_),
    .X(_2032_));
 sky130_fd_sc_hd__a21oi_2 _5277_ (.A1(_1777_),
    .A2(_2024_),
    .B1(_2032_),
    .Y(_2033_));
 sky130_fd_sc_hd__or2_2 _5278_ (.A(_1639_),
    .B(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__and2_2 _5279_ (.A(_1799_),
    .B(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__or2_2 _5280_ (.A(_2017_),
    .B(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__mux2_2 _5281_ (.A0(_1999_),
    .A1(_2036_),
    .S(_1877_),
    .X(_2037_));
 sky130_fd_sc_hd__mux2_2 _5282_ (.A0(_1962_),
    .A1(_2037_),
    .S(_1879_),
    .X(_2038_));
 sky130_fd_sc_hd__a32oi_2 _5283_ (.A1(_1171_),
    .A2(_1094_),
    .A3(_1098_),
    .B1(_1102_),
    .B2(_1109_),
    .Y(_2039_));
 sky130_fd_sc_hd__buf_1 _5284_ (.A(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__mux2_2 _5285_ (.A0(_1880_),
    .A1(_2038_),
    .S(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__mux4_2 _5286_ (.A0(\rf.registers[20][3] ),
    .A1(\rf.registers[21][3] ),
    .A2(\rf.registers[22][3] ),
    .A3(\rf.registers[23][3] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2042_));
 sky130_fd_sc_hd__mux4_2 _5287_ (.A0(\rf.registers[16][3] ),
    .A1(\rf.registers[17][3] ),
    .A2(\rf.registers[18][3] ),
    .A3(\rf.registers[19][3] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2043_));
 sky130_fd_sc_hd__buf_1 _5288_ (.A(_1684_),
    .X(_2044_));
 sky130_fd_sc_hd__mux2_2 _5289_ (.A0(_2042_),
    .A1(_2043_),
    .S(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__mux4_2 _5290_ (.A0(\rf.registers[28][3] ),
    .A1(\rf.registers[29][3] ),
    .A2(\rf.registers[30][3] ),
    .A3(\rf.registers[31][3] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2046_));
 sky130_fd_sc_hd__mux4_2 _5291_ (.A0(\rf.registers[24][3] ),
    .A1(\rf.registers[25][3] ),
    .A2(\rf.registers[26][3] ),
    .A3(\rf.registers[27][3] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2047_));
 sky130_fd_sc_hd__mux2_2 _5292_ (.A0(_2046_),
    .A1(_2047_),
    .S(_2044_),
    .X(_2048_));
 sky130_fd_sc_hd__mux2_2 _5293_ (.A0(_2045_),
    .A1(_2048_),
    .S(_1696_),
    .X(_2049_));
 sky130_fd_sc_hd__buf_1 _5294_ (.A(_1673_),
    .X(_2050_));
 sky130_fd_sc_hd__buf_1 _5295_ (.A(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__buf_1 _5296_ (.A(_1690_),
    .X(_2052_));
 sky130_fd_sc_hd__buf_1 _5297_ (.A(_2052_),
    .X(_2053_));
 sky130_fd_sc_hd__mux4_2 _5298_ (.A0(\rf.registers[8][3] ),
    .A1(\rf.registers[9][3] ),
    .A2(\rf.registers[10][3] ),
    .A3(\rf.registers[11][3] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__mux4_2 _5299_ (.A0(\rf.registers[12][3] ),
    .A1(\rf.registers[13][3] ),
    .A2(\rf.registers[14][3] ),
    .A3(\rf.registers[15][3] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2055_));
 sky130_fd_sc_hd__mux2_2 _5300_ (.A0(_2054_),
    .A1(_2055_),
    .S(_1712_),
    .X(_2056_));
 sky130_fd_sc_hd__nor2_2 _5301_ (.A(_1828_),
    .B(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__mux4_2 _5302_ (.A0(\rf.registers[4][3] ),
    .A1(\rf.registers[5][3] ),
    .A2(\rf.registers[6][3] ),
    .A3(\rf.registers[7][3] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2058_));
 sky130_fd_sc_hd__mux4_2 _5303_ (.A0(\rf.registers[0][3] ),
    .A1(\rf.registers[1][3] ),
    .A2(\rf.registers[2][3] ),
    .A3(\rf.registers[3][3] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2059_));
 sky130_fd_sc_hd__mux2_2 _5304_ (.A0(_2058_),
    .A1(_2059_),
    .S(_1685_),
    .X(_2060_));
 sky130_fd_sc_hd__o21ai_2 _5305_ (.A1(_1699_),
    .A2(_2060_),
    .B1(_1670_),
    .Y(_2061_));
 sky130_fd_sc_hd__o2bb2a_2 _5306_ (.A1_N(_1729_),
    .A2_N(_2049_),
    .B1(_2057_),
    .B2(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__or2_2 _5307_ (.A(_1638_),
    .B(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__or2_2 _5308_ (.A(_1167_),
    .B(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__mux4_2 _5309_ (.A0(\rf.registers[20][2] ),
    .A1(\rf.registers[21][2] ),
    .A2(\rf.registers[22][2] ),
    .A3(\rf.registers[23][2] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2065_));
 sky130_fd_sc_hd__mux4_2 _5310_ (.A0(\rf.registers[16][2] ),
    .A1(\rf.registers[17][2] ),
    .A2(\rf.registers[18][2] ),
    .A3(\rf.registers[19][2] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2066_));
 sky130_fd_sc_hd__mux2_2 _5311_ (.A0(_2065_),
    .A1(_2066_),
    .S(_1645_),
    .X(_2067_));
 sky130_fd_sc_hd__mux4_2 _5312_ (.A0(\rf.registers[28][2] ),
    .A1(\rf.registers[29][2] ),
    .A2(\rf.registers[30][2] ),
    .A3(\rf.registers[31][2] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2068_));
 sky130_fd_sc_hd__mux4_2 _5313_ (.A0(\rf.registers[24][2] ),
    .A1(\rf.registers[25][2] ),
    .A2(\rf.registers[26][2] ),
    .A3(\rf.registers[27][2] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2069_));
 sky130_fd_sc_hd__mux2_2 _5314_ (.A0(_2068_),
    .A1(_2069_),
    .S(_1645_),
    .X(_2070_));
 sky130_fd_sc_hd__mux2_2 _5315_ (.A0(_2067_),
    .A1(_2070_),
    .S(A1[3]),
    .X(_2071_));
 sky130_fd_sc_hd__mux4_2 _5316_ (.A0(\rf.registers[8][2] ),
    .A1(\rf.registers[9][2] ),
    .A2(\rf.registers[10][2] ),
    .A3(\rf.registers[11][2] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2072_));
 sky130_fd_sc_hd__and2_2 _5317_ (.A(_1684_),
    .B(_2072_),
    .X(_2073_));
 sky130_fd_sc_hd__mux4_2 _5318_ (.A0(\rf.registers[12][2] ),
    .A1(\rf.registers[13][2] ),
    .A2(\rf.registers[14][2] ),
    .A3(\rf.registers[15][2] ),
    .S0(_1673_),
    .S1(_1690_),
    .X(_2074_));
 sky130_fd_sc_hd__a21o_2 _5319_ (.A1(A1[2]),
    .A2(_2074_),
    .B1(_1655_),
    .X(_2075_));
 sky130_fd_sc_hd__mux4_2 _5320_ (.A0(\rf.registers[4][2] ),
    .A1(\rf.registers[5][2] ),
    .A2(\rf.registers[6][2] ),
    .A3(\rf.registers[7][2] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2076_));
 sky130_fd_sc_hd__mux4_2 _5321_ (.A0(\rf.registers[0][2] ),
    .A1(\rf.registers[1][2] ),
    .A2(\rf.registers[2][2] ),
    .A3(\rf.registers[3][2] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2077_));
 sky130_fd_sc_hd__mux2_2 _5322_ (.A0(_2076_),
    .A1(_2077_),
    .S(_1684_),
    .X(_2078_));
 sky130_fd_sc_hd__o221a_2 _5323_ (.A1(_2073_),
    .A2(_2075_),
    .B1(_2078_),
    .B2(A1[3]),
    .C1(_1640_),
    .X(_2079_));
 sky130_fd_sc_hd__a21oi_2 _5324_ (.A1(A1[4]),
    .A2(_2071_),
    .B1(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__nor2_2 _5325_ (.A(_1638_),
    .B(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2_2 _5326_ (.A(_1168_),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__and2_2 _5327_ (.A(_2064_),
    .B(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__mux4_2 _5328_ (.A0(\rf.registers[24][1] ),
    .A1(\rf.registers[25][1] ),
    .A2(\rf.registers[26][1] ),
    .A3(\rf.registers[27][1] ),
    .S0(_1673_),
    .S1(_1690_),
    .X(_2084_));
 sky130_fd_sc_hd__mux4_2 _5329_ (.A0(\rf.registers[28][1] ),
    .A1(\rf.registers[29][1] ),
    .A2(\rf.registers[30][1] ),
    .A3(\rf.registers[31][1] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2085_));
 sky130_fd_sc_hd__mux4_2 _5330_ (.A0(\rf.registers[16][1] ),
    .A1(\rf.registers[17][1] ),
    .A2(\rf.registers[18][1] ),
    .A3(\rf.registers[19][1] ),
    .S0(_1673_),
    .S1(_1690_),
    .X(_2086_));
 sky130_fd_sc_hd__mux4_2 _5331_ (.A0(\rf.registers[20][1] ),
    .A1(\rf.registers[21][1] ),
    .A2(\rf.registers[22][1] ),
    .A3(\rf.registers[23][1] ),
    .S0(_1673_),
    .S1(_1690_),
    .X(_2087_));
 sky130_fd_sc_hd__mux4_2 _5332_ (.A0(_2084_),
    .A1(_2085_),
    .A2(_2086_),
    .A3(_2087_),
    .S0(A1[2]),
    .S1(_1655_),
    .X(_2088_));
 sky130_fd_sc_hd__mux4_2 _5333_ (.A0(\rf.registers[4][1] ),
    .A1(\rf.registers[5][1] ),
    .A2(\rf.registers[6][1] ),
    .A3(\rf.registers[7][1] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_2089_));
 sky130_fd_sc_hd__or2_2 _5334_ (.A(_1645_),
    .B(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__mux4_2 _5335_ (.A0(\rf.registers[0][1] ),
    .A1(\rf.registers[1][1] ),
    .A2(\rf.registers[2][1] ),
    .A3(\rf.registers[3][1] ),
    .S0(_1701_),
    .S1(_1677_),
    .X(_2091_));
 sky130_fd_sc_hd__o21a_2 _5336_ (.A1(A1[2]),
    .A2(_2091_),
    .B1(_1655_),
    .X(_2092_));
 sky130_fd_sc_hd__mux4_2 _5337_ (.A0(\rf.registers[8][1] ),
    .A1(\rf.registers[9][1] ),
    .A2(\rf.registers[10][1] ),
    .A3(\rf.registers[11][1] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_2093_));
 sky130_fd_sc_hd__mux4_2 _5338_ (.A0(\rf.registers[12][1] ),
    .A1(\rf.registers[13][1] ),
    .A2(\rf.registers[14][1] ),
    .A3(\rf.registers[15][1] ),
    .S0(_1641_),
    .S1(_1642_),
    .X(_2094_));
 sky130_fd_sc_hd__mux2_2 _5339_ (.A0(_2093_),
    .A1(_2094_),
    .S(A1[2]),
    .X(_2095_));
 sky130_fd_sc_hd__a221o_2 _5340_ (.A1(_2090_),
    .A2(_2092_),
    .B1(_2095_),
    .B2(A1[3]),
    .C1(A1[4]),
    .X(_2096_));
 sky130_fd_sc_hd__o21ai_2 _5341_ (.A1(_1640_),
    .A2(_2088_),
    .B1(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__or2_2 _5342_ (.A(_1638_),
    .B(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__or2_2 _5343_ (.A(_1167_),
    .B(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__mux2_2 _5344_ (.A0(_2083_),
    .A1(_2099_),
    .S(_1148_),
    .X(_2100_));
 sky130_fd_sc_hd__nor2_2 _5345_ (.A(_1664_),
    .B(_1084_),
    .Y(_2101_));
 sky130_fd_sc_hd__nand2_2 _5346_ (.A(_1060_),
    .B(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__a31o_2 _5347_ (.A1(_1127_),
    .A2(_1663_),
    .A3(_2100_),
    .B1(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__buf_1 _5348_ (.A(_1111_),
    .X(_2104_));
 sky130_fd_sc_hd__buf_1 _5349_ (.A(_2104_),
    .X(_2105_));
 sky130_fd_sc_hd__mux4_2 _5350_ (.A0(\rf.registers[20][15] ),
    .A1(\rf.registers[21][15] ),
    .A2(\rf.registers[22][15] ),
    .A3(\rf.registers[23][15] ),
    .S0(_1734_),
    .S1(_1680_),
    .X(_2106_));
 sky130_fd_sc_hd__mux4_2 _5351_ (.A0(\rf.registers[16][15] ),
    .A1(\rf.registers[17][15] ),
    .A2(\rf.registers[18][15] ),
    .A3(\rf.registers[19][15] ),
    .S0(_1782_),
    .S1(_1680_),
    .X(_2107_));
 sky130_fd_sc_hd__mux4_2 _5352_ (.A0(\rf.registers[28][15] ),
    .A1(\rf.registers[29][15] ),
    .A2(\rf.registers[30][15] ),
    .A3(\rf.registers[31][15] ),
    .S0(_1782_),
    .S1(_1680_),
    .X(_2108_));
 sky130_fd_sc_hd__mux4_2 _5353_ (.A0(\rf.registers[24][15] ),
    .A1(\rf.registers[25][15] ),
    .A2(\rf.registers[26][15] ),
    .A3(\rf.registers[27][15] ),
    .S0(_1782_),
    .S1(_1680_),
    .X(_2109_));
 sky130_fd_sc_hd__mux4_2 _5354_ (.A0(_2106_),
    .A1(_2107_),
    .A2(_2108_),
    .A3(_2109_),
    .S0(_1685_),
    .S1(_1696_),
    .X(_2110_));
 sky130_fd_sc_hd__mux4_2 _5355_ (.A0(\rf.registers[8][15] ),
    .A1(\rf.registers[9][15] ),
    .A2(\rf.registers[10][15] ),
    .A3(\rf.registers[11][15] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2111_));
 sky130_fd_sc_hd__or2_2 _5356_ (.A(_1712_),
    .B(_2111_),
    .X(_2112_));
 sky130_fd_sc_hd__buf_1 _5357_ (.A(_1702_),
    .X(_2113_));
 sky130_fd_sc_hd__buf_1 _5358_ (.A(_2052_),
    .X(_2114_));
 sky130_fd_sc_hd__mux4_2 _5359_ (.A0(\rf.registers[12][15] ),
    .A1(\rf.registers[13][15] ),
    .A2(\rf.registers[14][15] ),
    .A3(\rf.registers[15][15] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__o21a_2 _5360_ (.A1(_1685_),
    .A2(_2115_),
    .B1(_1696_),
    .X(_2116_));
 sky130_fd_sc_hd__buf_1 _5361_ (.A(_1702_),
    .X(_2117_));
 sky130_fd_sc_hd__buf_1 _5362_ (.A(_1678_),
    .X(_2118_));
 sky130_fd_sc_hd__mux4_2 _5363_ (.A0(\rf.registers[4][15] ),
    .A1(\rf.registers[5][15] ),
    .A2(\rf.registers[6][15] ),
    .A3(\rf.registers[7][15] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__mux4_2 _5364_ (.A0(\rf.registers[0][15] ),
    .A1(\rf.registers[1][15] ),
    .A2(\rf.registers[2][15] ),
    .A3(\rf.registers[3][15] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2120_));
 sky130_fd_sc_hd__mux2_2 _5365_ (.A0(_2119_),
    .A1(_2120_),
    .S(_1738_),
    .X(_2121_));
 sky130_fd_sc_hd__a221o_2 _5366_ (.A1(_2112_),
    .A2(_2116_),
    .B1(_2121_),
    .B2(_1828_),
    .C1(_1728_),
    .X(_2122_));
 sky130_fd_sc_hd__o21ai_2 _5367_ (.A1(_1671_),
    .A2(_2110_),
    .B1(_2122_),
    .Y(_2123_));
 sky130_fd_sc_hd__nor2_2 _5368_ (.A(_1639_),
    .B(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__mux4_2 _5369_ (.A0(\rf.registers[20][14] ),
    .A1(\rf.registers[21][14] ),
    .A2(\rf.registers[22][14] ),
    .A3(\rf.registers[23][14] ),
    .S0(_1733_),
    .S1(_1679_),
    .X(_2125_));
 sky130_fd_sc_hd__mux4_2 _5370_ (.A0(\rf.registers[16][14] ),
    .A1(\rf.registers[17][14] ),
    .A2(\rf.registers[18][14] ),
    .A3(\rf.registers[19][14] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2126_));
 sky130_fd_sc_hd__mux2_2 _5371_ (.A0(_2125_),
    .A1(_2126_),
    .S(_2044_),
    .X(_2127_));
 sky130_fd_sc_hd__mux4_2 _5372_ (.A0(\rf.registers[28][14] ),
    .A1(\rf.registers[29][14] ),
    .A2(\rf.registers[30][14] ),
    .A3(\rf.registers[31][14] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2128_));
 sky130_fd_sc_hd__mux4_2 _5373_ (.A0(\rf.registers[24][14] ),
    .A1(\rf.registers[25][14] ),
    .A2(\rf.registers[26][14] ),
    .A3(\rf.registers[27][14] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2129_));
 sky130_fd_sc_hd__mux2_2 _5374_ (.A0(_2128_),
    .A1(_2129_),
    .S(_2044_),
    .X(_2130_));
 sky130_fd_sc_hd__mux2_2 _5375_ (.A0(_2127_),
    .A1(_2130_),
    .S(_1696_),
    .X(_2131_));
 sky130_fd_sc_hd__mux4_2 _5376_ (.A0(\rf.registers[8][14] ),
    .A1(\rf.registers[9][14] ),
    .A2(\rf.registers[10][14] ),
    .A3(\rf.registers[11][14] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2132_));
 sky130_fd_sc_hd__mux4_2 _5377_ (.A0(\rf.registers[12][14] ),
    .A1(\rf.registers[13][14] ),
    .A2(\rf.registers[14][14] ),
    .A3(\rf.registers[15][14] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2133_));
 sky130_fd_sc_hd__mux2_2 _5378_ (.A0(_2132_),
    .A1(_2133_),
    .S(_1711_),
    .X(_2134_));
 sky130_fd_sc_hd__nand2_2 _5379_ (.A(_1699_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__mux4_2 _5380_ (.A0(\rf.registers[4][14] ),
    .A1(\rf.registers[5][14] ),
    .A2(\rf.registers[6][14] ),
    .A3(\rf.registers[7][14] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2136_));
 sky130_fd_sc_hd__mux4_2 _5381_ (.A0(\rf.registers[0][14] ),
    .A1(\rf.registers[1][14] ),
    .A2(\rf.registers[2][14] ),
    .A3(\rf.registers[3][14] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2137_));
 sky130_fd_sc_hd__mux2_2 _5382_ (.A0(_2136_),
    .A1(_2137_),
    .S(_1738_),
    .X(_2138_));
 sky130_fd_sc_hd__a21oi_2 _5383_ (.A1(_1828_),
    .A2(_2138_),
    .B1(_1728_),
    .Y(_2139_));
 sky130_fd_sc_hd__a2bb2o_2 _5384_ (.A1_N(_1670_),
    .A2_N(_2131_),
    .B1(_2135_),
    .B2(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__nor2_2 _5385_ (.A(_1639_),
    .B(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__nor2_2 _5386_ (.A(_1669_),
    .B(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__o21ba_2 _5387_ (.A1(_1169_),
    .A2(_2124_),
    .B1_N(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__inv_2 _5388_ (.A(_1638_),
    .Y(_2144_));
 sky130_fd_sc_hd__mux4_2 _5389_ (.A0(\rf.registers[20][13] ),
    .A1(\rf.registers[21][13] ),
    .A2(\rf.registers[22][13] ),
    .A3(\rf.registers[23][13] ),
    .S0(_1673_),
    .S1(_1690_),
    .X(_2145_));
 sky130_fd_sc_hd__mux4_2 _5390_ (.A0(\rf.registers[16][13] ),
    .A1(\rf.registers[17][13] ),
    .A2(\rf.registers[18][13] ),
    .A3(\rf.registers[19][13] ),
    .S0(_1673_),
    .S1(_1690_),
    .X(_2146_));
 sky130_fd_sc_hd__mux2_2 _5391_ (.A0(_2145_),
    .A1(_2146_),
    .S(_1684_),
    .X(_2147_));
 sky130_fd_sc_hd__mux4_2 _5392_ (.A0(\rf.registers[28][13] ),
    .A1(\rf.registers[29][13] ),
    .A2(\rf.registers[30][13] ),
    .A3(\rf.registers[31][13] ),
    .S0(_1673_),
    .S1(_1690_),
    .X(_2148_));
 sky130_fd_sc_hd__mux4_2 _5393_ (.A0(\rf.registers[24][13] ),
    .A1(\rf.registers[25][13] ),
    .A2(\rf.registers[26][13] ),
    .A3(\rf.registers[27][13] ),
    .S0(_1673_),
    .S1(_1690_),
    .X(_2149_));
 sky130_fd_sc_hd__mux2_2 _5394_ (.A0(_2148_),
    .A1(_2149_),
    .S(_1684_),
    .X(_2150_));
 sky130_fd_sc_hd__mux2_2 _5395_ (.A0(_2147_),
    .A1(_2150_),
    .S(A1[3]),
    .X(_2151_));
 sky130_fd_sc_hd__mux4_2 _5396_ (.A0(\rf.registers[4][13] ),
    .A1(\rf.registers[5][13] ),
    .A2(\rf.registers[6][13] ),
    .A3(\rf.registers[7][13] ),
    .S0(_1702_),
    .S1(_1678_),
    .X(_2152_));
 sky130_fd_sc_hd__or2_2 _5397_ (.A(_1684_),
    .B(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__mux4_2 _5398_ (.A0(\rf.registers[0][13] ),
    .A1(\rf.registers[1][13] ),
    .A2(\rf.registers[2][13] ),
    .A3(\rf.registers[3][13] ),
    .S0(_1702_),
    .S1(_1678_),
    .X(_2154_));
 sky130_fd_sc_hd__o21a_2 _5399_ (.A1(_1711_),
    .A2(_2154_),
    .B1(_1655_),
    .X(_2155_));
 sky130_fd_sc_hd__mux4_2 _5400_ (.A0(\rf.registers[8][13] ),
    .A1(\rf.registers[9][13] ),
    .A2(\rf.registers[10][13] ),
    .A3(\rf.registers[11][13] ),
    .S0(_1702_),
    .S1(_1678_),
    .X(_2156_));
 sky130_fd_sc_hd__mux4_2 _5401_ (.A0(\rf.registers[12][13] ),
    .A1(\rf.registers[13][13] ),
    .A2(\rf.registers[14][13] ),
    .A3(\rf.registers[15][13] ),
    .S0(_1702_),
    .S1(_1678_),
    .X(_2157_));
 sky130_fd_sc_hd__mux2_2 _5402_ (.A0(_2156_),
    .A1(_2157_),
    .S(A1[2]),
    .X(_2158_));
 sky130_fd_sc_hd__a221o_2 _5403_ (.A1(_2153_),
    .A2(_2155_),
    .B1(_2158_),
    .B2(A1[3]),
    .C1(A1[4]),
    .X(_2159_));
 sky130_fd_sc_hd__o21a_2 _5404_ (.A1(_1640_),
    .A2(_2151_),
    .B1(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__a21oi_2 _5405_ (.A1(_2144_),
    .A2(_2160_),
    .B1(_1800_),
    .Y(_2161_));
 sky130_fd_sc_hd__mux4_2 _5406_ (.A0(\rf.registers[24][12] ),
    .A1(\rf.registers[25][12] ),
    .A2(\rf.registers[26][12] ),
    .A3(\rf.registers[27][12] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2162_));
 sky130_fd_sc_hd__mux4_2 _5407_ (.A0(\rf.registers[28][12] ),
    .A1(\rf.registers[29][12] ),
    .A2(\rf.registers[30][12] ),
    .A3(\rf.registers[31][12] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2163_));
 sky130_fd_sc_hd__mux4_2 _5408_ (.A0(\rf.registers[16][12] ),
    .A1(\rf.registers[17][12] ),
    .A2(\rf.registers[18][12] ),
    .A3(\rf.registers[19][12] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2164_));
 sky130_fd_sc_hd__mux4_2 _5409_ (.A0(\rf.registers[20][12] ),
    .A1(\rf.registers[21][12] ),
    .A2(\rf.registers[22][12] ),
    .A3(\rf.registers[23][12] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2165_));
 sky130_fd_sc_hd__mux4_2 _5410_ (.A0(_2162_),
    .A1(_2163_),
    .A2(_2164_),
    .A3(_2165_),
    .S0(_1711_),
    .S1(_1716_),
    .X(_2166_));
 sky130_fd_sc_hd__mux4_2 _5411_ (.A0(\rf.registers[8][12] ),
    .A1(\rf.registers[9][12] ),
    .A2(\rf.registers[10][12] ),
    .A3(\rf.registers[11][12] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2167_));
 sky130_fd_sc_hd__mux4_2 _5412_ (.A0(\rf.registers[12][12] ),
    .A1(\rf.registers[13][12] ),
    .A2(\rf.registers[14][12] ),
    .A3(\rf.registers[15][12] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2168_));
 sky130_fd_sc_hd__mux2_2 _5413_ (.A0(_2167_),
    .A1(_2168_),
    .S(_1711_),
    .X(_2169_));
 sky130_fd_sc_hd__nand2_2 _5414_ (.A(_1699_),
    .B(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__mux4_2 _5415_ (.A0(\rf.registers[4][12] ),
    .A1(\rf.registers[5][12] ),
    .A2(\rf.registers[6][12] ),
    .A3(\rf.registers[7][12] ),
    .S0(_1718_),
    .S1(_1721_),
    .X(_2171_));
 sky130_fd_sc_hd__mux4_2 _5416_ (.A0(\rf.registers[0][12] ),
    .A1(\rf.registers[1][12] ),
    .A2(\rf.registers[2][12] ),
    .A3(\rf.registers[3][12] ),
    .S0(_1718_),
    .S1(_1721_),
    .X(_2172_));
 sky130_fd_sc_hd__mux2_2 _5417_ (.A0(_2171_),
    .A1(_2172_),
    .S(_1738_),
    .X(_2173_));
 sky130_fd_sc_hd__a21oi_2 _5418_ (.A1(_1828_),
    .A2(_2173_),
    .B1(_1728_),
    .Y(_2174_));
 sky130_fd_sc_hd__a2bb2o_2 _5419_ (.A1_N(_1670_),
    .A2_N(_2166_),
    .B1(_2170_),
    .B2(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__o21ai_2 _5420_ (.A1(_1758_),
    .A2(_2175_),
    .B1(_1800_),
    .Y(_2176_));
 sky130_fd_sc_hd__and2b_2 _5421_ (.A_N(_2161_),
    .B(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__buf_1 _5422_ (.A(_1877_),
    .X(_2178_));
 sky130_fd_sc_hd__mux2_2 _5423_ (.A0(_2143_),
    .A1(_2177_),
    .S(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__mux4_2 _5424_ (.A0(\rf.registers[24][11] ),
    .A1(\rf.registers[25][11] ),
    .A2(\rf.registers[26][11] ),
    .A3(\rf.registers[27][11] ),
    .S0(_1675_),
    .S1(_1692_),
    .X(_2180_));
 sky130_fd_sc_hd__mux4_2 _5425_ (.A0(\rf.registers[28][11] ),
    .A1(\rf.registers[29][11] ),
    .A2(\rf.registers[30][11] ),
    .A3(\rf.registers[31][11] ),
    .S0(_1675_),
    .S1(_1692_),
    .X(_2181_));
 sky130_fd_sc_hd__mux4_2 _5426_ (.A0(\rf.registers[16][11] ),
    .A1(\rf.registers[17][11] ),
    .A2(\rf.registers[18][11] ),
    .A3(\rf.registers[19][11] ),
    .S0(_1675_),
    .S1(_1692_),
    .X(_2182_));
 sky130_fd_sc_hd__mux4_2 _5427_ (.A0(\rf.registers[20][11] ),
    .A1(\rf.registers[21][11] ),
    .A2(\rf.registers[22][11] ),
    .A3(\rf.registers[23][11] ),
    .S0(_1675_),
    .S1(_1692_),
    .X(_2183_));
 sky130_fd_sc_hd__mux4_2 _5428_ (.A0(_2180_),
    .A1(_2181_),
    .A2(_2182_),
    .A3(_2183_),
    .S0(_1712_),
    .S1(_1716_),
    .X(_2184_));
 sky130_fd_sc_hd__mux4_2 _5429_ (.A0(\rf.registers[12][11] ),
    .A1(\rf.registers[13][11] ),
    .A2(\rf.registers[14][11] ),
    .A3(\rf.registers[15][11] ),
    .S0(_1704_),
    .S1(_1707_),
    .X(_2185_));
 sky130_fd_sc_hd__mux4_2 _5430_ (.A0(\rf.registers[8][11] ),
    .A1(\rf.registers[9][11] ),
    .A2(\rf.registers[10][11] ),
    .A3(\rf.registers[11][11] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2186_));
 sky130_fd_sc_hd__or2_2 _5431_ (.A(_1711_),
    .B(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__o211a_2 _5432_ (.A1(_1686_),
    .A2(_2185_),
    .B1(_2187_),
    .C1(_1699_),
    .X(_2188_));
 sky130_fd_sc_hd__mux4_2 _5433_ (.A0(\rf.registers[4][11] ),
    .A1(\rf.registers[5][11] ),
    .A2(\rf.registers[6][11] ),
    .A3(\rf.registers[7][11] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2189_));
 sky130_fd_sc_hd__mux4_2 _5434_ (.A0(\rf.registers[0][11] ),
    .A1(\rf.registers[1][11] ),
    .A2(\rf.registers[2][11] ),
    .A3(\rf.registers[3][11] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2190_));
 sky130_fd_sc_hd__mux2_2 _5435_ (.A0(_2189_),
    .A1(_2190_),
    .S(_1738_),
    .X(_2191_));
 sky130_fd_sc_hd__a21o_2 _5436_ (.A1(_1828_),
    .A2(_2191_),
    .B1(_1728_),
    .X(_2192_));
 sky130_fd_sc_hd__o22a_2 _5437_ (.A1(_1670_),
    .A2(_2184_),
    .B1(_2188_),
    .B2(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__and2_2 _5438_ (.A(_2144_),
    .B(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__mux4_2 _5439_ (.A0(\rf.registers[24][10] ),
    .A1(\rf.registers[25][10] ),
    .A2(\rf.registers[26][10] ),
    .A3(\rf.registers[27][10] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2195_));
 sky130_fd_sc_hd__mux4_2 _5440_ (.A0(\rf.registers[28][10] ),
    .A1(\rf.registers[29][10] ),
    .A2(\rf.registers[30][10] ),
    .A3(\rf.registers[31][10] ),
    .S0(_1674_),
    .S1(_1691_),
    .X(_2196_));
 sky130_fd_sc_hd__mux2_2 _5441_ (.A0(_2195_),
    .A1(_2196_),
    .S(_1711_),
    .X(_2197_));
 sky130_fd_sc_hd__mux4_2 _5442_ (.A0(\rf.registers[20][10] ),
    .A1(\rf.registers[21][10] ),
    .A2(\rf.registers[22][10] ),
    .A3(\rf.registers[23][10] ),
    .S0(_2050_),
    .S1(_2052_),
    .X(_2198_));
 sky130_fd_sc_hd__mux4_2 _5443_ (.A0(\rf.registers[16][10] ),
    .A1(\rf.registers[17][10] ),
    .A2(\rf.registers[18][10] ),
    .A3(\rf.registers[19][10] ),
    .S0(_2050_),
    .S1(_2052_),
    .X(_2199_));
 sky130_fd_sc_hd__mux2_2 _5444_ (.A0(_2198_),
    .A1(_2199_),
    .S(_2044_),
    .X(_2200_));
 sky130_fd_sc_hd__mux2_2 _5445_ (.A0(_2197_),
    .A1(_2200_),
    .S(_1716_),
    .X(_2201_));
 sky130_fd_sc_hd__mux4_2 _5446_ (.A0(\rf.registers[8][10] ),
    .A1(\rf.registers[9][10] ),
    .A2(\rf.registers[10][10] ),
    .A3(\rf.registers[11][10] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2202_));
 sky130_fd_sc_hd__mux4_2 _5447_ (.A0(\rf.registers[12][10] ),
    .A1(\rf.registers[13][10] ),
    .A2(\rf.registers[14][10] ),
    .A3(\rf.registers[15][10] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2203_));
 sky130_fd_sc_hd__mux2_2 _5448_ (.A0(_2202_),
    .A1(_2203_),
    .S(_1711_),
    .X(_2204_));
 sky130_fd_sc_hd__nand2_2 _5449_ (.A(_1699_),
    .B(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__mux4_2 _5450_ (.A0(\rf.registers[4][10] ),
    .A1(\rf.registers[5][10] ),
    .A2(\rf.registers[6][10] ),
    .A3(\rf.registers[7][10] ),
    .S0(_1718_),
    .S1(_1721_),
    .X(_2206_));
 sky130_fd_sc_hd__mux4_2 _5451_ (.A0(\rf.registers[0][10] ),
    .A1(\rf.registers[1][10] ),
    .A2(\rf.registers[2][10] ),
    .A3(\rf.registers[3][10] ),
    .S0(_1718_),
    .S1(_1721_),
    .X(_2207_));
 sky130_fd_sc_hd__mux2_2 _5452_ (.A0(_2206_),
    .A1(_2207_),
    .S(_1738_),
    .X(_2208_));
 sky130_fd_sc_hd__a21oi_2 _5453_ (.A1(_1828_),
    .A2(_2208_),
    .B1(_1728_),
    .Y(_2209_));
 sky130_fd_sc_hd__a2bb2o_2 _5454_ (.A1_N(_1670_),
    .A2_N(_2201_),
    .B1(_2205_),
    .B2(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__or2_2 _5455_ (.A(_1639_),
    .B(_2210_),
    .X(_2211_));
 sky130_fd_sc_hd__and2_2 _5456_ (.A(_1168_),
    .B(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__o21ba_2 _5457_ (.A1(_1169_),
    .A2(_2194_),
    .B1_N(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__mux4_2 _5458_ (.A0(\rf.registers[20][8] ),
    .A1(\rf.registers[21][8] ),
    .A2(\rf.registers[22][8] ),
    .A3(\rf.registers[23][8] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2214_));
 sky130_fd_sc_hd__mux4_2 _5459_ (.A0(\rf.registers[16][8] ),
    .A1(\rf.registers[17][8] ),
    .A2(\rf.registers[18][8] ),
    .A3(\rf.registers[19][8] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2215_));
 sky130_fd_sc_hd__mux2_2 _5460_ (.A0(_2214_),
    .A1(_2215_),
    .S(_1685_),
    .X(_2216_));
 sky130_fd_sc_hd__mux4_2 _5461_ (.A0(\rf.registers[28][8] ),
    .A1(\rf.registers[29][8] ),
    .A2(\rf.registers[30][8] ),
    .A3(\rf.registers[31][8] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2217_));
 sky130_fd_sc_hd__mux4_2 _5462_ (.A0(\rf.registers[24][8] ),
    .A1(\rf.registers[25][8] ),
    .A2(\rf.registers[26][8] ),
    .A3(\rf.registers[27][8] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2218_));
 sky130_fd_sc_hd__mux2_2 _5463_ (.A0(_2217_),
    .A1(_2218_),
    .S(_1685_),
    .X(_2219_));
 sky130_fd_sc_hd__mux2_2 _5464_ (.A0(_2216_),
    .A1(_2219_),
    .S(_1699_),
    .X(_2220_));
 sky130_fd_sc_hd__mux4_2 _5465_ (.A0(\rf.registers[8][8] ),
    .A1(\rf.registers[9][8] ),
    .A2(\rf.registers[10][8] ),
    .A3(\rf.registers[11][8] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_2221_));
 sky130_fd_sc_hd__mux4_2 _5466_ (.A0(\rf.registers[12][8] ),
    .A1(\rf.registers[13][8] ),
    .A2(\rf.registers[14][8] ),
    .A3(\rf.registers[15][8] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_2222_));
 sky130_fd_sc_hd__mux2_2 _5467_ (.A0(_2221_),
    .A1(_2222_),
    .S(_1712_),
    .X(_2223_));
 sky130_fd_sc_hd__nand2_2 _5468_ (.A(_1697_),
    .B(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hd__mux4_2 _5469_ (.A0(\rf.registers[4][8] ),
    .A1(\rf.registers[5][8] ),
    .A2(\rf.registers[6][8] ),
    .A3(\rf.registers[7][8] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_2225_));
 sky130_fd_sc_hd__mux4_2 _5470_ (.A0(\rf.registers[0][8] ),
    .A1(\rf.registers[1][8] ),
    .A2(\rf.registers[2][8] ),
    .A3(\rf.registers[3][8] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_2226_));
 sky130_fd_sc_hd__mux2_2 _5471_ (.A0(_2225_),
    .A1(_2226_),
    .S(_1739_),
    .X(_2227_));
 sky130_fd_sc_hd__a21oi_2 _5472_ (.A1(_1717_),
    .A2(_2227_),
    .B1(_1729_),
    .Y(_2228_));
 sky130_fd_sc_hd__a2bb2o_2 _5473_ (.A1_N(_1671_),
    .A2_N(_2220_),
    .B1(_2224_),
    .B2(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__or2_2 _5474_ (.A(_1639_),
    .B(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__mux4_2 _5475_ (.A0(\rf.registers[24][9] ),
    .A1(\rf.registers[25][9] ),
    .A2(\rf.registers[26][9] ),
    .A3(\rf.registers[27][9] ),
    .S0(_1675_),
    .S1(_1692_),
    .X(_2231_));
 sky130_fd_sc_hd__mux4_2 _5476_ (.A0(\rf.registers[28][9] ),
    .A1(\rf.registers[29][9] ),
    .A2(\rf.registers[30][9] ),
    .A3(\rf.registers[31][9] ),
    .S0(_1675_),
    .S1(_1692_),
    .X(_2232_));
 sky130_fd_sc_hd__mux2_2 _5477_ (.A0(_2231_),
    .A1(_2232_),
    .S(_1712_),
    .X(_2233_));
 sky130_fd_sc_hd__mux4_2 _5478_ (.A0(\rf.registers[20][9] ),
    .A1(\rf.registers[21][9] ),
    .A2(\rf.registers[22][9] ),
    .A3(\rf.registers[23][9] ),
    .S0(_1675_),
    .S1(_1692_),
    .X(_2234_));
 sky130_fd_sc_hd__mux4_2 _5479_ (.A0(\rf.registers[16][9] ),
    .A1(\rf.registers[17][9] ),
    .A2(\rf.registers[18][9] ),
    .A3(\rf.registers[19][9] ),
    .S0(_1675_),
    .S1(_1692_),
    .X(_2235_));
 sky130_fd_sc_hd__mux2_2 _5480_ (.A0(_2234_),
    .A1(_2235_),
    .S(_1685_),
    .X(_2236_));
 sky130_fd_sc_hd__mux2_2 _5481_ (.A0(_2233_),
    .A1(_2236_),
    .S(_1828_),
    .X(_2237_));
 sky130_fd_sc_hd__mux4_2 _5482_ (.A0(\rf.registers[12][9] ),
    .A1(\rf.registers[13][9] ),
    .A2(\rf.registers[14][9] ),
    .A3(\rf.registers[15][9] ),
    .S0(_1782_),
    .S1(_1680_),
    .X(_2238_));
 sky130_fd_sc_hd__mux4_2 _5483_ (.A0(\rf.registers[8][9] ),
    .A1(\rf.registers[9][9] ),
    .A2(\rf.registers[10][9] ),
    .A3(\rf.registers[11][9] ),
    .S0(_1782_),
    .S1(_1692_),
    .X(_2239_));
 sky130_fd_sc_hd__mux2_2 _5484_ (.A0(_2238_),
    .A1(_2239_),
    .S(_1685_),
    .X(_2240_));
 sky130_fd_sc_hd__mux4_2 _5485_ (.A0(\rf.registers[4][9] ),
    .A1(\rf.registers[5][9] ),
    .A2(\rf.registers[6][9] ),
    .A3(\rf.registers[7][9] ),
    .S0(_1734_),
    .S1(_1735_),
    .X(_2241_));
 sky130_fd_sc_hd__or2_2 _5486_ (.A(_1739_),
    .B(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__mux4_2 _5487_ (.A0(\rf.registers[0][9] ),
    .A1(\rf.registers[1][9] ),
    .A2(\rf.registers[2][9] ),
    .A3(\rf.registers[3][9] ),
    .S0(_1719_),
    .S1(_1722_),
    .X(_2243_));
 sky130_fd_sc_hd__o21a_2 _5488_ (.A1(_1712_),
    .A2(_2243_),
    .B1(_1716_),
    .X(_2244_));
 sky130_fd_sc_hd__a221o_2 _5489_ (.A1(_1697_),
    .A2(_2240_),
    .B1(_2242_),
    .B2(_2244_),
    .C1(_1729_),
    .X(_2245_));
 sky130_fd_sc_hd__o21ai_2 _5490_ (.A1(_1671_),
    .A2(_2237_),
    .B1(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__nor2_2 _5491_ (.A(_1842_),
    .B(_2246_),
    .Y(_2247_));
 sky130_fd_sc_hd__nand2_2 _5492_ (.A(_1668_),
    .B(_2247_),
    .Y(_2248_));
 sky130_fd_sc_hd__o21ai_2 _5493_ (.A1(_1669_),
    .A2(_2230_),
    .B1(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__mux2_2 _5494_ (.A0(_2213_),
    .A1(_2249_),
    .S(_2178_),
    .X(_2250_));
 sky130_fd_sc_hd__buf_1 _5495_ (.A(_1125_),
    .X(_2251_));
 sky130_fd_sc_hd__buf_1 _5496_ (.A(_2251_),
    .X(_2252_));
 sky130_fd_sc_hd__mux2_2 _5497_ (.A0(_2179_),
    .A1(_2250_),
    .S(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__or2_2 _5498_ (.A(_2039_),
    .B(_1126_),
    .X(_2254_));
 sky130_fd_sc_hd__buf_1 _5499_ (.A(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__mux4_2 _5500_ (.A0(\rf.registers[20][6] ),
    .A1(\rf.registers[21][6] ),
    .A2(\rf.registers[22][6] ),
    .A3(\rf.registers[23][6] ),
    .S0(_1733_),
    .S1(_1679_),
    .X(_2256_));
 sky130_fd_sc_hd__mux4_2 _5501_ (.A0(\rf.registers[16][6] ),
    .A1(\rf.registers[17][6] ),
    .A2(\rf.registers[18][6] ),
    .A3(\rf.registers[19][6] ),
    .S0(_1733_),
    .S1(_1679_),
    .X(_2257_));
 sky130_fd_sc_hd__mux2_2 _5502_ (.A0(_2256_),
    .A1(_2257_),
    .S(_2044_),
    .X(_2258_));
 sky130_fd_sc_hd__mux4_2 _5503_ (.A0(\rf.registers[28][6] ),
    .A1(\rf.registers[29][6] ),
    .A2(\rf.registers[30][6] ),
    .A3(\rf.registers[31][6] ),
    .S0(_1733_),
    .S1(_1679_),
    .X(_2259_));
 sky130_fd_sc_hd__mux4_2 _5504_ (.A0(\rf.registers[24][6] ),
    .A1(\rf.registers[25][6] ),
    .A2(\rf.registers[26][6] ),
    .A3(\rf.registers[27][6] ),
    .S0(_1733_),
    .S1(_1679_),
    .X(_2260_));
 sky130_fd_sc_hd__mux2_2 _5505_ (.A0(_2259_),
    .A1(_2260_),
    .S(_2044_),
    .X(_2261_));
 sky130_fd_sc_hd__mux2_2 _5506_ (.A0(_2258_),
    .A1(_2261_),
    .S(_1696_),
    .X(_2262_));
 sky130_fd_sc_hd__mux4_2 _5507_ (.A0(\rf.registers[8][6] ),
    .A1(\rf.registers[9][6] ),
    .A2(\rf.registers[10][6] ),
    .A3(\rf.registers[11][6] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2263_));
 sky130_fd_sc_hd__mux4_2 _5508_ (.A0(\rf.registers[12][6] ),
    .A1(\rf.registers[13][6] ),
    .A2(\rf.registers[14][6] ),
    .A3(\rf.registers[15][6] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2264_));
 sky130_fd_sc_hd__mux2_2 _5509_ (.A0(_2263_),
    .A1(_2264_),
    .S(_1712_),
    .X(_2265_));
 sky130_fd_sc_hd__nand2_2 _5510_ (.A(_1699_),
    .B(_2265_),
    .Y(_2266_));
 sky130_fd_sc_hd__mux4_2 _5511_ (.A0(\rf.registers[4][6] ),
    .A1(\rf.registers[5][6] ),
    .A2(\rf.registers[6][6] ),
    .A3(\rf.registers[7][6] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2267_));
 sky130_fd_sc_hd__mux4_2 _5512_ (.A0(\rf.registers[0][6] ),
    .A1(\rf.registers[1][6] ),
    .A2(\rf.registers[2][6] ),
    .A3(\rf.registers[3][6] ),
    .S0(_1703_),
    .S1(_1706_),
    .X(_2268_));
 sky130_fd_sc_hd__mux2_2 _5513_ (.A0(_2267_),
    .A1(_2268_),
    .S(_1738_),
    .X(_2269_));
 sky130_fd_sc_hd__a21oi_2 _5514_ (.A1(_1828_),
    .A2(_2269_),
    .B1(_1728_),
    .Y(_2270_));
 sky130_fd_sc_hd__a2bb2o_2 _5515_ (.A1_N(_1670_),
    .A2_N(_2262_),
    .B1(_2266_),
    .B2(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__or2_2 _5516_ (.A(_1638_),
    .B(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__mux4_2 _5517_ (.A0(\rf.registers[24][7] ),
    .A1(\rf.registers[25][7] ),
    .A2(\rf.registers[26][7] ),
    .A3(\rf.registers[27][7] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2273_));
 sky130_fd_sc_hd__mux4_2 _5518_ (.A0(\rf.registers[28][7] ),
    .A1(\rf.registers[29][7] ),
    .A2(\rf.registers[30][7] ),
    .A3(\rf.registers[31][7] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2274_));
 sky130_fd_sc_hd__mux4_2 _5519_ (.A0(\rf.registers[16][7] ),
    .A1(\rf.registers[17][7] ),
    .A2(\rf.registers[18][7] ),
    .A3(\rf.registers[19][7] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2275_));
 sky130_fd_sc_hd__mux4_2 _5520_ (.A0(\rf.registers[20][7] ),
    .A1(\rf.registers[21][7] ),
    .A2(\rf.registers[22][7] ),
    .A3(\rf.registers[23][7] ),
    .S0(_2051_),
    .S1(_2053_),
    .X(_2276_));
 sky130_fd_sc_hd__mux4_2 _5521_ (.A0(_2273_),
    .A1(_2274_),
    .A2(_2275_),
    .A3(_2276_),
    .S0(_1711_),
    .S1(_1716_),
    .X(_2277_));
 sky130_fd_sc_hd__mux4_2 _5522_ (.A0(\rf.registers[12][7] ),
    .A1(\rf.registers[13][7] ),
    .A2(\rf.registers[14][7] ),
    .A3(\rf.registers[15][7] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2278_));
 sky130_fd_sc_hd__mux4_2 _5523_ (.A0(\rf.registers[8][7] ),
    .A1(\rf.registers[9][7] ),
    .A2(\rf.registers[10][7] ),
    .A3(\rf.registers[11][7] ),
    .S0(_2113_),
    .S1(_2114_),
    .X(_2279_));
 sky130_fd_sc_hd__mux2_2 _5524_ (.A0(_2278_),
    .A1(_2279_),
    .S(_1685_),
    .X(_2280_));
 sky130_fd_sc_hd__nand2_2 _5525_ (.A(_1699_),
    .B(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__mux4_2 _5526_ (.A0(\rf.registers[4][7] ),
    .A1(\rf.registers[5][7] ),
    .A2(\rf.registers[6][7] ),
    .A3(\rf.registers[7][7] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2282_));
 sky130_fd_sc_hd__mux4_2 _5527_ (.A0(\rf.registers[0][7] ),
    .A1(\rf.registers[1][7] ),
    .A2(\rf.registers[2][7] ),
    .A3(\rf.registers[3][7] ),
    .S0(_2117_),
    .S1(_2118_),
    .X(_2283_));
 sky130_fd_sc_hd__mux2_2 _5528_ (.A0(_2282_),
    .A1(_2283_),
    .S(_1738_),
    .X(_2284_));
 sky130_fd_sc_hd__a21oi_2 _5529_ (.A1(_1828_),
    .A2(_2284_),
    .B1(_1728_),
    .Y(_2285_));
 sky130_fd_sc_hd__a2bb2o_2 _5530_ (.A1_N(_1670_),
    .A2_N(_2277_),
    .B1(_2281_),
    .B2(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__nor2_2 _5531_ (.A(_1638_),
    .B(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__nor2_2 _5532_ (.A(_1800_),
    .B(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__a21oi_2 _5533_ (.A1(_1169_),
    .A2(_2272_),
    .B1(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__mux4_2 _5534_ (.A0(\rf.registers[20][4] ),
    .A1(\rf.registers[21][4] ),
    .A2(\rf.registers[22][4] ),
    .A3(\rf.registers[23][4] ),
    .S0(_2050_),
    .S1(_2052_),
    .X(_2290_));
 sky130_fd_sc_hd__mux4_2 _5535_ (.A0(\rf.registers[16][4] ),
    .A1(\rf.registers[17][4] ),
    .A2(\rf.registers[18][4] ),
    .A3(\rf.registers[19][4] ),
    .S0(_2050_),
    .S1(_2052_),
    .X(_2291_));
 sky130_fd_sc_hd__mux2_2 _5536_ (.A0(_2290_),
    .A1(_2291_),
    .S(_2044_),
    .X(_2292_));
 sky130_fd_sc_hd__mux4_2 _5537_ (.A0(\rf.registers[28][4] ),
    .A1(\rf.registers[29][4] ),
    .A2(\rf.registers[30][4] ),
    .A3(\rf.registers[31][4] ),
    .S0(_2050_),
    .S1(_2052_),
    .X(_2293_));
 sky130_fd_sc_hd__mux4_2 _5538_ (.A0(\rf.registers[24][4] ),
    .A1(\rf.registers[25][4] ),
    .A2(\rf.registers[26][4] ),
    .A3(\rf.registers[27][4] ),
    .S0(_2050_),
    .S1(_2052_),
    .X(_2294_));
 sky130_fd_sc_hd__mux2_2 _5539_ (.A0(_2293_),
    .A1(_2294_),
    .S(_2044_),
    .X(_2295_));
 sky130_fd_sc_hd__mux2_2 _5540_ (.A0(_2292_),
    .A1(_2295_),
    .S(_1696_),
    .X(_2296_));
 sky130_fd_sc_hd__mux4_2 _5541_ (.A0(\rf.registers[12][4] ),
    .A1(\rf.registers[13][4] ),
    .A2(\rf.registers[14][4] ),
    .A3(\rf.registers[15][4] ),
    .S0(_1718_),
    .S1(_1721_),
    .X(_2297_));
 sky130_fd_sc_hd__mux4_2 _5542_ (.A0(\rf.registers[8][4] ),
    .A1(\rf.registers[9][4] ),
    .A2(\rf.registers[10][4] ),
    .A3(\rf.registers[11][4] ),
    .S0(_1718_),
    .S1(_1721_),
    .X(_2298_));
 sky130_fd_sc_hd__mux2_2 _5543_ (.A0(_2297_),
    .A1(_2298_),
    .S(_1738_),
    .X(_2299_));
 sky130_fd_sc_hd__nor2_2 _5544_ (.A(_1716_),
    .B(_2299_),
    .Y(_2300_));
 sky130_fd_sc_hd__mux4_2 _5545_ (.A0(\rf.registers[4][4] ),
    .A1(\rf.registers[5][4] ),
    .A2(\rf.registers[6][4] ),
    .A3(\rf.registers[7][4] ),
    .S0(_1718_),
    .S1(_1679_),
    .X(_2301_));
 sky130_fd_sc_hd__mux4_2 _5546_ (.A0(\rf.registers[0][4] ),
    .A1(\rf.registers[1][4] ),
    .A2(\rf.registers[2][4] ),
    .A3(\rf.registers[3][4] ),
    .S0(_1733_),
    .S1(_1679_),
    .X(_2302_));
 sky130_fd_sc_hd__mux2_2 _5547_ (.A0(_2301_),
    .A1(_2302_),
    .S(_1738_),
    .X(_2303_));
 sky130_fd_sc_hd__o21ai_2 _5548_ (.A1(_1696_),
    .A2(_2303_),
    .B1(_1670_),
    .Y(_2304_));
 sky130_fd_sc_hd__o2bb2a_2 _5549_ (.A1_N(_1728_),
    .A2_N(_2296_),
    .B1(_2300_),
    .B2(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__nor2_2 _5550_ (.A(_1842_),
    .B(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__nand2_2 _5551_ (.A(_1799_),
    .B(_2306_),
    .Y(_2307_));
 sky130_fd_sc_hd__mux4_2 _5552_ (.A0(\rf.registers[20][5] ),
    .A1(\rf.registers[21][5] ),
    .A2(\rf.registers[22][5] ),
    .A3(\rf.registers[23][5] ),
    .S0(_2050_),
    .S1(_2052_),
    .X(_2308_));
 sky130_fd_sc_hd__mux4_2 _5553_ (.A0(\rf.registers[16][5] ),
    .A1(\rf.registers[17][5] ),
    .A2(\rf.registers[18][5] ),
    .A3(\rf.registers[19][5] ),
    .S0(_2050_),
    .S1(_2052_),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_2 _5554_ (.A0(_2308_),
    .A1(_2309_),
    .S(_1684_),
    .X(_2310_));
 sky130_fd_sc_hd__mux4_2 _5555_ (.A0(\rf.registers[28][5] ),
    .A1(\rf.registers[29][5] ),
    .A2(\rf.registers[30][5] ),
    .A3(\rf.registers[31][5] ),
    .S0(_2050_),
    .S1(_1678_),
    .X(_2311_));
 sky130_fd_sc_hd__mux4_2 _5556_ (.A0(\rf.registers[24][5] ),
    .A1(\rf.registers[25][5] ),
    .A2(\rf.registers[26][5] ),
    .A3(\rf.registers[27][5] ),
    .S0(_1702_),
    .S1(_1678_),
    .X(_2312_));
 sky130_fd_sc_hd__mux2_2 _5557_ (.A0(_2311_),
    .A1(_2312_),
    .S(_1684_),
    .X(_2313_));
 sky130_fd_sc_hd__mux2_2 _5558_ (.A0(_2310_),
    .A1(_2313_),
    .S(A1[3]),
    .X(_2314_));
 sky130_fd_sc_hd__mux4_2 _5559_ (.A0(\rf.registers[8][5] ),
    .A1(\rf.registers[9][5] ),
    .A2(\rf.registers[10][5] ),
    .A3(\rf.registers[11][5] ),
    .S0(_1718_),
    .S1(_1721_),
    .X(_2315_));
 sky130_fd_sc_hd__mux4_2 _5560_ (.A0(\rf.registers[12][5] ),
    .A1(\rf.registers[13][5] ),
    .A2(\rf.registers[14][5] ),
    .A3(\rf.registers[15][5] ),
    .S0(_1718_),
    .S1(_1721_),
    .X(_2316_));
 sky130_fd_sc_hd__mux2_2 _5561_ (.A0(_2315_),
    .A1(_2316_),
    .S(_1711_),
    .X(_2317_));
 sky130_fd_sc_hd__nor2_2 _5562_ (.A(_1716_),
    .B(_2317_),
    .Y(_2318_));
 sky130_fd_sc_hd__mux4_2 _5563_ (.A0(\rf.registers[4][5] ),
    .A1(\rf.registers[5][5] ),
    .A2(\rf.registers[6][5] ),
    .A3(\rf.registers[7][5] ),
    .S0(_1733_),
    .S1(_1679_),
    .X(_2319_));
 sky130_fd_sc_hd__mux4_2 _5564_ (.A0(\rf.registers[0][5] ),
    .A1(\rf.registers[1][5] ),
    .A2(\rf.registers[2][5] ),
    .A3(\rf.registers[3][5] ),
    .S0(_1733_),
    .S1(_1679_),
    .X(_2320_));
 sky130_fd_sc_hd__mux2_2 _5565_ (.A0(_2319_),
    .A1(_2320_),
    .S(_2044_),
    .X(_2321_));
 sky130_fd_sc_hd__o21ai_2 _5566_ (.A1(_1696_),
    .A2(_2321_),
    .B1(_1670_),
    .Y(_2322_));
 sky130_fd_sc_hd__o2bb2a_2 _5567_ (.A1_N(_1728_),
    .A2_N(_2314_),
    .B1(_2318_),
    .B2(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__nor2_2 _5568_ (.A(_1842_),
    .B(_2323_),
    .Y(_2324_));
 sky130_fd_sc_hd__nand2_2 _5569_ (.A(_1839_),
    .B(_2324_),
    .Y(_2325_));
 sky130_fd_sc_hd__nand2_2 _5570_ (.A(_2307_),
    .B(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__buf_1 _5571_ (.A(_1803_),
    .X(_2327_));
 sky130_fd_sc_hd__mux2_2 _5572_ (.A0(_2289_),
    .A1(_2326_),
    .S(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__o22ai_2 _5573_ (.A1(_2105_),
    .A2(_2253_),
    .B1(_2255_),
    .B2(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__o22a_2 _5574_ (.A1(_1666_),
    .A2(_2041_),
    .B1(_2103_),
    .B2(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__or2_2 _5575_ (.A(_1669_),
    .B(_1660_),
    .X(_2331_));
 sky130_fd_sc_hd__nand2_2 _5576_ (.A(_1669_),
    .B(_1660_),
    .Y(_2332_));
 sky130_fd_sc_hd__buf_1 _5577_ (.A(opcode[1]),
    .X(_2333_));
 sky130_fd_sc_hd__a21o_2 _5578_ (.A1(_2331_),
    .A2(_2332_),
    .B1(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__o211ai_2 _5579_ (.A1(_1128_),
    .A2(_1663_),
    .B1(_2330_),
    .C1(_2334_),
    .Y(alu_out[0]));
 sky130_fd_sc_hd__nand2_2 _5580_ (.A(_1060_),
    .B(_1085_),
    .Y(_2335_));
 sky130_fd_sc_hd__nand2_2 _5581_ (.A(_1111_),
    .B(_1126_),
    .Y(_2336_));
 sky130_fd_sc_hd__buf_1 _5582_ (.A(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__nor2_2 _5583_ (.A(_1167_),
    .B(_1661_),
    .Y(_2338_));
 sky130_fd_sc_hd__a21oi_2 _5584_ (.A1(_1799_),
    .A2(_2098_),
    .B1(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__nand2_2 _5585_ (.A(_2178_),
    .B(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__o21a_2 _5586_ (.A1(_1758_),
    .A2(_1874_),
    .B1(_1839_),
    .X(_2341_));
 sky130_fd_sc_hd__or2_2 _5587_ (.A(_1667_),
    .B(_2124_),
    .X(_2342_));
 sky130_fd_sc_hd__and2b_2 _5588_ (.A_N(_2341_),
    .B(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__or2_2 _5589_ (.A(_1799_),
    .B(_2141_),
    .X(_2344_));
 sky130_fd_sc_hd__a21o_2 _5590_ (.A1(_2144_),
    .A2(_2160_),
    .B1(_1668_),
    .X(_2345_));
 sky130_fd_sc_hd__and2_2 _5591_ (.A(_2344_),
    .B(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__buf_1 _5592_ (.A(_1146_),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_2 _5593_ (.A0(_2343_),
    .A1(_2346_),
    .S(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__o21ai_2 _5594_ (.A1(_1758_),
    .A2(_2175_),
    .B1(_1839_),
    .Y(_2349_));
 sky130_fd_sc_hd__or2_2 _5595_ (.A(_1668_),
    .B(_2194_),
    .X(_2350_));
 sky130_fd_sc_hd__and2_2 _5596_ (.A(_2349_),
    .B(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__nand2_2 _5597_ (.A(_1839_),
    .B(_2211_),
    .Y(_2352_));
 sky130_fd_sc_hd__or2_2 _5598_ (.A(_1668_),
    .B(_2247_),
    .X(_2353_));
 sky130_fd_sc_hd__and2_2 _5599_ (.A(_2352_),
    .B(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__mux2_2 _5600_ (.A0(_2351_),
    .A1(_2354_),
    .S(_2347_),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_2 _5601_ (.A0(_2348_),
    .A1(_2355_),
    .S(_1879_),
    .X(_2356_));
 sky130_fd_sc_hd__or2_2 _5602_ (.A(_1667_),
    .B(_2287_),
    .X(_2357_));
 sky130_fd_sc_hd__nand2_2 _5603_ (.A(_1839_),
    .B(_2230_),
    .Y(_2358_));
 sky130_fd_sc_hd__and2_2 _5604_ (.A(_2357_),
    .B(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__or2_2 _5605_ (.A(_1668_),
    .B(_2324_),
    .X(_2360_));
 sky130_fd_sc_hd__nand2_2 _5606_ (.A(_1667_),
    .B(_2272_),
    .Y(_2361_));
 sky130_fd_sc_hd__and2_2 _5607_ (.A(_2360_),
    .B(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__buf_1 _5608_ (.A(_1877_),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_2 _5609_ (.A0(_2359_),
    .A1(_2362_),
    .S(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__a21bo_2 _5610_ (.A1(_1169_),
    .A2(_2098_),
    .B1_N(_1803_),
    .X(_2365_));
 sky130_fd_sc_hd__inv_2 _5611_ (.A(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__or2_2 _5612_ (.A(_1167_),
    .B(_2081_),
    .X(_2367_));
 sky130_fd_sc_hd__nand2_2 _5613_ (.A(_1167_),
    .B(_2063_),
    .Y(_2368_));
 sky130_fd_sc_hd__or2_2 _5614_ (.A(_1799_),
    .B(_2306_),
    .X(_2369_));
 sky130_fd_sc_hd__and3b_2 _5615_ (.A_N(_2363_),
    .B(_2368_),
    .C(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__a211o_2 _5616_ (.A1(_2366_),
    .A2(_2367_),
    .B1(_2370_),
    .C1(_2336_),
    .X(_2371_));
 sky130_fd_sc_hd__and2_2 _5617_ (.A(_1060_),
    .B(_2101_),
    .X(_2372_));
 sky130_fd_sc_hd__buf_1 _5618_ (.A(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__o211a_2 _5619_ (.A1(_2255_),
    .A2(_2364_),
    .B1(_2371_),
    .C1(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__o21ai_2 _5620_ (.A1(_2105_),
    .A2(_2356_),
    .B1(_2374_),
    .Y(_2375_));
 sky130_fd_sc_hd__o311a_2 _5621_ (.A1(_2335_),
    .A2(_2337_),
    .A3(_2340_),
    .B1(_2375_),
    .C1(_2333_),
    .X(_2376_));
 sky130_fd_sc_hd__and2_2 _5622_ (.A(_1168_),
    .B(_1905_),
    .X(_2377_));
 sky130_fd_sc_hd__inv_2 _5623_ (.A(_2377_),
    .Y(_2378_));
 sky130_fd_sc_hd__nor2_2 _5624_ (.A(_1799_),
    .B(_1924_),
    .Y(_2379_));
 sky130_fd_sc_hd__and2_2 _5625_ (.A(_1167_),
    .B(_1943_),
    .X(_2380_));
 sky130_fd_sc_hd__nor2_2 _5626_ (.A(_2379_),
    .B(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__mux2_2 _5627_ (.A0(_2378_),
    .A1(_2381_),
    .S(_1877_),
    .X(_2382_));
 sky130_fd_sc_hd__nand2_2 _5628_ (.A(_1668_),
    .B(_1959_),
    .Y(_2383_));
 sky130_fd_sc_hd__nand2_2 _5629_ (.A(_1799_),
    .B(_1979_),
    .Y(_2384_));
 sky130_fd_sc_hd__nand2_2 _5630_ (.A(_2383_),
    .B(_2384_),
    .Y(_2385_));
 sky130_fd_sc_hd__and2_2 _5631_ (.A(_1167_),
    .B(_2016_),
    .X(_2386_));
 sky130_fd_sc_hd__o21ba_2 _5632_ (.A1(_1168_),
    .A2(_1997_),
    .B1_N(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_2 _5633_ (.A0(_2385_),
    .A1(_2387_),
    .S(_1145_),
    .X(_2388_));
 sky130_fd_sc_hd__inv_2 _5634_ (.A(_2388_),
    .Y(_2389_));
 sky130_fd_sc_hd__mux2_2 _5635_ (.A0(_2382_),
    .A1(_2389_),
    .S(_2251_),
    .X(_2390_));
 sky130_fd_sc_hd__and2_2 _5636_ (.A(_1667_),
    .B(_2034_),
    .X(_2391_));
 sky130_fd_sc_hd__and2_2 _5637_ (.A(_1799_),
    .B(_1732_),
    .X(_2392_));
 sky130_fd_sc_hd__nor2_2 _5638_ (.A(_2391_),
    .B(_2392_),
    .Y(_2393_));
 sky130_fd_sc_hd__nor2_2 _5639_ (.A(_1168_),
    .B(_1755_),
    .Y(_2394_));
 sky130_fd_sc_hd__nor2_2 _5640_ (.A(_1668_),
    .B(_1780_),
    .Y(_2395_));
 sky130_fd_sc_hd__nor2_2 _5641_ (.A(_2394_),
    .B(_2395_),
    .Y(_2396_));
 sky130_fd_sc_hd__mux2_2 _5642_ (.A0(_2393_),
    .A1(_2396_),
    .S(_1146_),
    .X(_2397_));
 sky130_fd_sc_hd__o21a_2 _5643_ (.A1(_1842_),
    .A2(_1798_),
    .B1(_1667_),
    .X(_2398_));
 sky130_fd_sc_hd__o21ai_2 _5644_ (.A1(_1842_),
    .A2(_1838_),
    .B1(_1799_),
    .Y(_2399_));
 sky130_fd_sc_hd__and2b_2 _5645_ (.A_N(_2398_),
    .B(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__nor2_2 _5646_ (.A(_1667_),
    .B(_1859_),
    .Y(_2401_));
 sky130_fd_sc_hd__o21ba_2 _5647_ (.A1(_1168_),
    .A2(_1821_),
    .B1_N(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__mux2_2 _5648_ (.A0(_2400_),
    .A1(_2402_),
    .S(_1145_),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_2 _5649_ (.A0(_2397_),
    .A1(_2403_),
    .S(_1125_),
    .X(_2404_));
 sky130_fd_sc_hd__inv_2 _5650_ (.A(_2404_),
    .Y(_2405_));
 sky130_fd_sc_hd__mux2_2 _5651_ (.A0(_2390_),
    .A1(_2405_),
    .S(_2104_),
    .X(_2406_));
 sky130_fd_sc_hd__or2_2 _5652_ (.A(_1666_),
    .B(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__buf_1 _5653_ (.A(_2333_),
    .X(_2408_));
 sky130_fd_sc_hd__nor2_2 _5654_ (.A(_1664_),
    .B(opcode[1]),
    .Y(_2409_));
 sky130_fd_sc_hd__or3_2 _5655_ (.A(_1145_),
    .B(_1166_),
    .C(_2409_),
    .X(_2410_));
 sky130_fd_sc_hd__buf_1 _5656_ (.A(_2409_),
    .X(_2411_));
 sky130_fd_sc_hd__o21ai_2 _5657_ (.A1(_1166_),
    .A2(_2411_),
    .B1(_1145_),
    .Y(_2412_));
 sky130_fd_sc_hd__a21oi_2 _5658_ (.A1(_2410_),
    .A2(_2412_),
    .B1(_2097_),
    .Y(_2413_));
 sky130_fd_sc_hd__and3_2 _5659_ (.A(_2097_),
    .B(_2410_),
    .C(_2412_),
    .X(_2414_));
 sky130_fd_sc_hd__or2_2 _5660_ (.A(_2413_),
    .B(_2414_),
    .X(_2415_));
 sky130_fd_sc_hd__xnor2_2 _5661_ (.A(_2332_),
    .B(_2415_),
    .Y(_2416_));
 sky130_fd_sc_hd__o2bb2a_2 _5662_ (.A1_N(_2376_),
    .A2_N(_2407_),
    .B1(_2408_),
    .B2(_2416_),
    .X(alu_out[1]));
 sky130_fd_sc_hd__inv_2 _5663_ (.A(_1662_),
    .Y(_2417_));
 sky130_fd_sc_hd__nand2_2 _5664_ (.A(_2082_),
    .B(_2099_),
    .Y(_2418_));
 sky130_fd_sc_hd__nand2_2 _5665_ (.A(_1147_),
    .B(_2418_),
    .Y(_2419_));
 sky130_fd_sc_hd__o21a_2 _5666_ (.A1(_2363_),
    .A2(_2417_),
    .B1(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__buf_1 _5667_ (.A(_2333_),
    .X(_2421_));
 sky130_fd_sc_hd__o21ai_2 _5668_ (.A1(_1128_),
    .A2(_2420_),
    .B1(_2421_),
    .Y(_2422_));
 sky130_fd_sc_hd__inv_2 _5669_ (.A(_1876_),
    .Y(_2423_));
 sky130_fd_sc_hd__mux2_2 _5670_ (.A0(_2423_),
    .A1(_2143_),
    .S(_1147_),
    .X(_2424_));
 sky130_fd_sc_hd__mux2_2 _5671_ (.A0(_2177_),
    .A1(_2213_),
    .S(_2363_),
    .X(_2425_));
 sky130_fd_sc_hd__buf_1 _5672_ (.A(_1879_),
    .X(_2426_));
 sky130_fd_sc_hd__mux2_2 _5673_ (.A0(_2424_),
    .A1(_2425_),
    .S(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__and2_2 _5674_ (.A(_1168_),
    .B(_2230_),
    .X(_2428_));
 sky130_fd_sc_hd__nor2_2 _5675_ (.A(_1800_),
    .B(_2247_),
    .Y(_2429_));
 sky130_fd_sc_hd__nor2_2 _5676_ (.A(_2428_),
    .B(_2429_),
    .Y(_2430_));
 sky130_fd_sc_hd__mux2_2 _5677_ (.A0(_2430_),
    .A1(_2289_),
    .S(_2363_),
    .X(_2431_));
 sky130_fd_sc_hd__inv_2 _5678_ (.A(_2083_),
    .Y(_2432_));
 sky130_fd_sc_hd__a21oi_2 _5679_ (.A1(_2307_),
    .A2(_2325_),
    .B1(_1148_),
    .Y(_2433_));
 sky130_fd_sc_hd__a211o_2 _5680_ (.A1(_1148_),
    .A2(_2432_),
    .B1(_2433_),
    .C1(_2337_),
    .X(_2434_));
 sky130_fd_sc_hd__o211a_2 _5681_ (.A1(_2255_),
    .A2(_2431_),
    .B1(_2434_),
    .C1(_2373_),
    .X(_2435_));
 sky130_fd_sc_hd__o21a_2 _5682_ (.A1(_2105_),
    .A2(_2427_),
    .B1(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__mux2_2 _5683_ (.A0(_2036_),
    .A1(_1757_),
    .S(_2347_),
    .X(_2437_));
 sky130_fd_sc_hd__or2b_2 _5684_ (.A(_1841_),
    .B_N(_2347_),
    .X(_2438_));
 sky130_fd_sc_hd__o21ai_2 _5685_ (.A1(_2178_),
    .A2(_1802_),
    .B1(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__nand2_2 _5686_ (.A(_2252_),
    .B(_2439_),
    .Y(_2440_));
 sky130_fd_sc_hd__o21a_2 _5687_ (.A1(_2252_),
    .A2(_2437_),
    .B1(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__or2b_2 _5688_ (.A(_1926_),
    .B_N(_2178_),
    .X(_2442_));
 sky130_fd_sc_hd__mux2_2 _5689_ (.A0(_1961_),
    .A1(_1999_),
    .S(_2347_),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_2 _5690_ (.A0(_2442_),
    .A1(_2443_),
    .S(_2252_),
    .X(_2444_));
 sky130_fd_sc_hd__mux2_2 _5691_ (.A0(_2441_),
    .A1(_2444_),
    .S(_2040_),
    .X(_2445_));
 sky130_fd_sc_hd__nor2_2 _5692_ (.A(_1666_),
    .B(_2445_),
    .Y(_2446_));
 sky130_fd_sc_hd__a21oi_2 _5693_ (.A1(_1145_),
    .A2(_1166_),
    .B1(_2411_),
    .Y(_2447_));
 sky130_fd_sc_hd__xnor2_2 _5694_ (.A(_1125_),
    .B(_2447_),
    .Y(_2448_));
 sky130_fd_sc_hd__xor2_2 _5695_ (.A(_2080_),
    .B(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__and2_2 _5696_ (.A(_1667_),
    .B(_1660_),
    .X(_2450_));
 sky130_fd_sc_hd__o21bai_2 _5697_ (.A1(_2450_),
    .A2(_2414_),
    .B1_N(_2413_),
    .Y(_2451_));
 sky130_fd_sc_hd__nand2_2 _5698_ (.A(_2449_),
    .B(_2451_),
    .Y(_2452_));
 sky130_fd_sc_hd__or2_2 _5699_ (.A(_2449_),
    .B(_2451_),
    .X(_2453_));
 sky130_fd_sc_hd__a21o_2 _5700_ (.A1(_2452_),
    .A2(_2453_),
    .B1(_2421_),
    .X(_2454_));
 sky130_fd_sc_hd__o31a_2 _5701_ (.A1(_2422_),
    .A2(_2436_),
    .A3(_2446_),
    .B1(_2454_),
    .X(alu_out[2]));
 sky130_fd_sc_hd__inv_2 _5702_ (.A(_2339_),
    .Y(_2455_));
 sky130_fd_sc_hd__and2_2 _5703_ (.A(_2368_),
    .B(_2367_),
    .X(_2456_));
 sky130_fd_sc_hd__inv_2 _5704_ (.A(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__mux2_2 _5705_ (.A0(_2455_),
    .A1(_2457_),
    .S(_1146_),
    .X(_2458_));
 sky130_fd_sc_hd__o21ai_2 _5706_ (.A1(_1128_),
    .A2(_2458_),
    .B1(_2421_),
    .Y(_2459_));
 sky130_fd_sc_hd__mux2_2 _5707_ (.A0(_2402_),
    .A1(_2343_),
    .S(_2327_),
    .X(_2460_));
 sky130_fd_sc_hd__mux2_2 _5708_ (.A0(_2346_),
    .A1(_2351_),
    .S(_2327_),
    .X(_2461_));
 sky130_fd_sc_hd__mux2_2 _5709_ (.A0(_2460_),
    .A1(_2461_),
    .S(_2252_),
    .X(_2462_));
 sky130_fd_sc_hd__mux2_2 _5710_ (.A0(_2354_),
    .A1(_2359_),
    .S(_2178_),
    .X(_2463_));
 sky130_fd_sc_hd__and2b_2 _5711_ (.A_N(_2178_),
    .B(_2362_),
    .X(_2464_));
 sky130_fd_sc_hd__a311o_2 _5712_ (.A1(_1148_),
    .A2(_2368_),
    .A3(_2369_),
    .B1(_2464_),
    .C1(_2336_),
    .X(_2465_));
 sky130_fd_sc_hd__o211a_2 _5713_ (.A1(_2255_),
    .A2(_2463_),
    .B1(_2465_),
    .C1(_2373_),
    .X(_2466_));
 sky130_fd_sc_hd__o21a_2 _5714_ (.A1(_2105_),
    .A2(_2462_),
    .B1(_2466_),
    .X(_2467_));
 sky130_fd_sc_hd__inv_2 _5715_ (.A(_1666_),
    .Y(_2468_));
 sky130_fd_sc_hd__mux2_2 _5716_ (.A0(_2387_),
    .A1(_2393_),
    .S(_1146_),
    .X(_2469_));
 sky130_fd_sc_hd__mux2_2 _5717_ (.A0(_2396_),
    .A1(_2400_),
    .S(_1877_),
    .X(_2470_));
 sky130_fd_sc_hd__mux2_2 _5718_ (.A0(_2469_),
    .A1(_2470_),
    .S(_2251_),
    .X(_2471_));
 sky130_fd_sc_hd__and3_2 _5719_ (.A(_2347_),
    .B(_1169_),
    .C(_1905_),
    .X(_2472_));
 sky130_fd_sc_hd__inv_2 _5720_ (.A(_2381_),
    .Y(_2473_));
 sky130_fd_sc_hd__mux2_2 _5721_ (.A0(_2473_),
    .A1(_2385_),
    .S(_1146_),
    .X(_2474_));
 sky130_fd_sc_hd__mux2_2 _5722_ (.A0(_2472_),
    .A1(_2474_),
    .S(_2251_),
    .X(_2475_));
 sky130_fd_sc_hd__mux2_2 _5723_ (.A0(_2471_),
    .A1(_2475_),
    .S(_2040_),
    .X(_2476_));
 sky130_fd_sc_hd__and2_2 _5724_ (.A(_2468_),
    .B(_2476_),
    .X(_2477_));
 sky130_fd_sc_hd__a31o_2 _5725_ (.A1(_1125_),
    .A2(_1145_),
    .A3(_1167_),
    .B1(_2411_),
    .X(_2478_));
 sky130_fd_sc_hd__xnor2_2 _5726_ (.A(_2039_),
    .B(_2478_),
    .Y(_2479_));
 sky130_fd_sc_hd__nor2_2 _5727_ (.A(_2062_),
    .B(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__nand2_2 _5728_ (.A(_2062_),
    .B(_2479_),
    .Y(_2481_));
 sky130_fd_sc_hd__or2b_2 _5729_ (.A(_2480_),
    .B_N(_2481_),
    .X(_2482_));
 sky130_fd_sc_hd__nor2_2 _5730_ (.A(_2080_),
    .B(_2448_),
    .Y(_2483_));
 sky130_fd_sc_hd__a21o_2 _5731_ (.A1(_2449_),
    .A2(_2451_),
    .B1(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__xnor2_2 _5732_ (.A(_2482_),
    .B(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hd__o32a_2 _5733_ (.A1(_2459_),
    .A2(_2467_),
    .A3(_2477_),
    .B1(_2485_),
    .B2(_2408_),
    .X(alu_out[3]));
 sky130_fd_sc_hd__mux2_2 _5734_ (.A0(_2037_),
    .A1(_1804_),
    .S(_2251_),
    .X(_2486_));
 sky130_fd_sc_hd__nand2_2 _5735_ (.A(_2039_),
    .B(_2251_),
    .Y(_2487_));
 sky130_fd_sc_hd__o22a_2 _5736_ (.A1(_2040_),
    .A2(_2486_),
    .B1(_2487_),
    .B2(_1962_),
    .X(_2488_));
 sky130_fd_sc_hd__nor2_2 _5737_ (.A(_1666_),
    .B(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__inv_2 _5738_ (.A(_1878_),
    .Y(_2490_));
 sky130_fd_sc_hd__mux2_2 _5739_ (.A0(_2490_),
    .A1(_2179_),
    .S(_2426_),
    .X(_2491_));
 sky130_fd_sc_hd__or2_2 _5740_ (.A(_2336_),
    .B(_2328_),
    .X(_2492_));
 sky130_fd_sc_hd__o211a_2 _5741_ (.A1(_2250_),
    .A2(_2255_),
    .B1(_2492_),
    .C1(_2373_),
    .X(_2493_));
 sky130_fd_sc_hd__o21a_2 _5742_ (.A1(_2105_),
    .A2(_2491_),
    .B1(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__nor2_2 _5743_ (.A(_2040_),
    .B(_2335_),
    .Y(_2495_));
 sky130_fd_sc_hd__buf_1 _5744_ (.A(_2495_),
    .X(_2496_));
 sky130_fd_sc_hd__and3_2 _5745_ (.A(_2327_),
    .B(_1169_),
    .C(_1661_),
    .X(_2497_));
 sky130_fd_sc_hd__and2_2 _5746_ (.A(_2064_),
    .B(_2307_),
    .X(_2498_));
 sky130_fd_sc_hd__inv_2 _5747_ (.A(_2498_),
    .Y(_2499_));
 sky130_fd_sc_hd__mux2_2 _5748_ (.A0(_2418_),
    .A1(_2499_),
    .S(_1147_),
    .X(_2500_));
 sky130_fd_sc_hd__buf_1 _5749_ (.A(_1126_),
    .X(_2501_));
 sky130_fd_sc_hd__mux2_2 _5750_ (.A0(_2497_),
    .A1(_2500_),
    .S(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__inv_2 _5751_ (.A(opcode[1]),
    .Y(_2503_));
 sky130_fd_sc_hd__buf_1 _5752_ (.A(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__a21o_2 _5753_ (.A1(_2496_),
    .A2(_2502_),
    .B1(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__and4_2 _5754_ (.A(_1110_),
    .B(_1125_),
    .C(_1144_),
    .D(_1166_),
    .X(_2506_));
 sky130_fd_sc_hd__nor2_2 _5755_ (.A(_2411_),
    .B(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__xnor2_2 _5756_ (.A(_1060_),
    .B(_2507_),
    .Y(_2508_));
 sky130_fd_sc_hd__nor2_2 _5757_ (.A(_2305_),
    .B(_2508_),
    .Y(_2509_));
 sky130_fd_sc_hd__and2_2 _5758_ (.A(_2305_),
    .B(_2508_),
    .X(_2510_));
 sky130_fd_sc_hd__nor2_2 _5759_ (.A(_2509_),
    .B(_2510_),
    .Y(_2511_));
 sky130_fd_sc_hd__a21o_2 _5760_ (.A1(_2481_),
    .A2(_2484_),
    .B1(_2480_),
    .X(_2512_));
 sky130_fd_sc_hd__xor2_2 _5761_ (.A(_2511_),
    .B(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__o32a_2 _5762_ (.A1(_2489_),
    .A2(_2494_),
    .A3(_2505_),
    .B1(_2513_),
    .B2(_2408_),
    .X(alu_out[4]));
 sky130_fd_sc_hd__a21oi_2 _5763_ (.A1(_1060_),
    .A2(_2506_),
    .B1(_2411_),
    .Y(_2514_));
 sky130_fd_sc_hd__xnor2_2 _5764_ (.A(_1083_),
    .B(_2514_),
    .Y(_2515_));
 sky130_fd_sc_hd__and2_2 _5765_ (.A(_2323_),
    .B(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__nor2_2 _5766_ (.A(_2323_),
    .B(_2515_),
    .Y(_2517_));
 sky130_fd_sc_hd__nor2_2 _5767_ (.A(_2516_),
    .B(_2517_),
    .Y(_2518_));
 sky130_fd_sc_hd__a21oi_2 _5768_ (.A1(_2511_),
    .A2(_2512_),
    .B1(_2509_),
    .Y(_2519_));
 sky130_fd_sc_hd__xnor2_2 _5769_ (.A(_2518_),
    .B(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__and2_2 _5770_ (.A(_2503_),
    .B(_2520_),
    .X(_2521_));
 sky130_fd_sc_hd__mux2_2 _5771_ (.A0(_2388_),
    .A1(_2397_),
    .S(_1126_),
    .X(_2522_));
 sky130_fd_sc_hd__o2bb2a_2 _5772_ (.A1_N(_1111_),
    .A2_N(_2522_),
    .B1(_2487_),
    .B2(_2382_),
    .X(_2523_));
 sky130_fd_sc_hd__nor2_2 _5773_ (.A(_2338_),
    .B(_2365_),
    .Y(_2524_));
 sky130_fd_sc_hd__nand2_2 _5774_ (.A(_2369_),
    .B(_2360_),
    .Y(_2525_));
 sky130_fd_sc_hd__nand2_2 _5775_ (.A(_2327_),
    .B(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__o21a_2 _5776_ (.A1(_2363_),
    .A2(_2456_),
    .B1(_2526_),
    .X(_2527_));
 sky130_fd_sc_hd__mux2_2 _5777_ (.A0(_2524_),
    .A1(_2527_),
    .S(_2501_),
    .X(_2528_));
 sky130_fd_sc_hd__a2bb2o_2 _5778_ (.A1_N(_1666_),
    .A2_N(_2523_),
    .B1(_2528_),
    .B2(_2495_),
    .X(_2529_));
 sky130_fd_sc_hd__buf_1 _5779_ (.A(_1111_),
    .X(_2530_));
 sky130_fd_sc_hd__mux2_2 _5780_ (.A0(_2403_),
    .A1(_2348_),
    .S(_1879_),
    .X(_2531_));
 sky130_fd_sc_hd__o22a_2 _5781_ (.A1(_2255_),
    .A2(_2355_),
    .B1(_2364_),
    .B2(_2337_),
    .X(_2532_));
 sky130_fd_sc_hd__o211a_2 _5782_ (.A1(_2530_),
    .A2(_2531_),
    .B1(_2532_),
    .C1(_2373_),
    .X(_2533_));
 sky130_fd_sc_hd__or3_2 _5783_ (.A(_2521_),
    .B(_2529_),
    .C(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__buf_1 _5784_ (.A(_2534_),
    .X(alu_out[5]));
 sky130_fd_sc_hd__and2_2 _5785_ (.A(_1059_),
    .B(_1083_),
    .X(_2535_));
 sky130_fd_sc_hd__buf_1 _5786_ (.A(_2411_),
    .X(_2536_));
 sky130_fd_sc_hd__a21oi_2 _5787_ (.A1(_2506_),
    .A2(_2535_),
    .B1(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__xnor2_2 _5788_ (.A(_1399_),
    .B(_2537_),
    .Y(_2538_));
 sky130_fd_sc_hd__and2_2 _5789_ (.A(_2271_),
    .B(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__nor2_2 _5790_ (.A(_2271_),
    .B(_2538_),
    .Y(_2540_));
 sky130_fd_sc_hd__nand2_2 _5791_ (.A(_2323_),
    .B(_2515_),
    .Y(_2541_));
 sky130_fd_sc_hd__a21o_2 _5792_ (.A1(_2509_),
    .A2(_2541_),
    .B1(_2517_),
    .X(_2542_));
 sky130_fd_sc_hd__a31oi_2 _5793_ (.A1(_2511_),
    .A2(_2512_),
    .A3(_2518_),
    .B1(_2542_),
    .Y(_2543_));
 sky130_fd_sc_hd__o21ai_2 _5794_ (.A1(_2539_),
    .A2(_2540_),
    .B1(_2543_),
    .Y(_2544_));
 sky130_fd_sc_hd__or3_2 _5795_ (.A(_2539_),
    .B(_2540_),
    .C(_2543_),
    .X(_2545_));
 sky130_fd_sc_hd__o31ai_2 _5796_ (.A1(_2363_),
    .A2(_1758_),
    .A3(_2331_),
    .B1(_2419_),
    .Y(_2546_));
 sky130_fd_sc_hd__o21ai_2 _5797_ (.A1(_1669_),
    .A2(_2272_),
    .B1(_2325_),
    .Y(_2547_));
 sky130_fd_sc_hd__mux2_2 _5798_ (.A0(_2499_),
    .A1(_2547_),
    .S(_2347_),
    .X(_2548_));
 sky130_fd_sc_hd__mux2_2 _5799_ (.A0(_2546_),
    .A1(_2548_),
    .S(_2501_),
    .X(_2549_));
 sky130_fd_sc_hd__mux2_2 _5800_ (.A0(_2439_),
    .A1(_2424_),
    .S(_2501_),
    .X(_2550_));
 sky130_fd_sc_hd__o22a_2 _5801_ (.A1(_2254_),
    .A2(_2425_),
    .B1(_2431_),
    .B2(_2337_),
    .X(_2551_));
 sky130_fd_sc_hd__o211a_2 _5802_ (.A1(_2530_),
    .A2(_2550_),
    .B1(_2551_),
    .C1(_2373_),
    .X(_2552_));
 sky130_fd_sc_hd__mux2_2 _5803_ (.A0(_2443_),
    .A1(_2437_),
    .S(_1879_),
    .X(_2553_));
 sky130_fd_sc_hd__o22a_2 _5804_ (.A1(_2442_),
    .A2(_2487_),
    .B1(_2553_),
    .B2(_2040_),
    .X(_2554_));
 sky130_fd_sc_hd__nor2_2 _5805_ (.A(_1666_),
    .B(_2554_),
    .Y(_2555_));
 sky130_fd_sc_hd__a211o_2 _5806_ (.A1(_2496_),
    .A2(_2549_),
    .B1(_2552_),
    .C1(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__a31o_2 _5807_ (.A1(_2504_),
    .A2(_2544_),
    .A3(_2545_),
    .B1(_2556_),
    .X(alu_out[6]));
 sky130_fd_sc_hd__a31o_2 _5808_ (.A1(_1399_),
    .A2(_2506_),
    .A3(_2535_),
    .B1(_2411_),
    .X(_2557_));
 sky130_fd_sc_hd__xor2_2 _5809_ (.A(_1415_),
    .B(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__and2_2 _5810_ (.A(_2286_),
    .B(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__or2_2 _5811_ (.A(_2286_),
    .B(_2558_),
    .X(_2560_));
 sky130_fd_sc_hd__or2b_2 _5812_ (.A(_2559_),
    .B_N(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__or2_2 _5813_ (.A(_2271_),
    .B(_2538_),
    .X(_2562_));
 sky130_fd_sc_hd__o21ai_2 _5814_ (.A1(_2539_),
    .A2(_2543_),
    .B1(_2562_),
    .Y(_2563_));
 sky130_fd_sc_hd__xnor2_2 _5815_ (.A(_2561_),
    .B(_2563_),
    .Y(_2564_));
 sky130_fd_sc_hd__and2_2 _5816_ (.A(_2361_),
    .B(_2357_),
    .X(_2565_));
 sky130_fd_sc_hd__inv_2 _5817_ (.A(_2565_),
    .Y(_2566_));
 sky130_fd_sc_hd__mux2_2 _5818_ (.A0(_2525_),
    .A1(_2566_),
    .S(_1146_),
    .X(_2567_));
 sky130_fd_sc_hd__mux2_2 _5819_ (.A0(_2458_),
    .A1(_2567_),
    .S(_1126_),
    .X(_2568_));
 sky130_fd_sc_hd__inv_2 _5820_ (.A(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__and2_2 _5821_ (.A(_2039_),
    .B(_2251_),
    .X(_2570_));
 sky130_fd_sc_hd__mux2_2 _5822_ (.A0(_2474_),
    .A1(_2469_),
    .S(_1126_),
    .X(_2571_));
 sky130_fd_sc_hd__a22o_2 _5823_ (.A1(_2472_),
    .A2(_2570_),
    .B1(_2571_),
    .B2(_1111_),
    .X(_2572_));
 sky130_fd_sc_hd__mux2_2 _5824_ (.A0(_2470_),
    .A1(_2460_),
    .S(_2252_),
    .X(_2573_));
 sky130_fd_sc_hd__o22a_2 _5825_ (.A1(_2255_),
    .A2(_2461_),
    .B1(_2463_),
    .B2(_2337_),
    .X(_2574_));
 sky130_fd_sc_hd__o211a_2 _5826_ (.A1(_2105_),
    .A2(_2573_),
    .B1(_2574_),
    .C1(_2373_),
    .X(_2575_));
 sky130_fd_sc_hd__a221o_2 _5827_ (.A1(_2496_),
    .A2(_2569_),
    .B1(_2572_),
    .B2(_2468_),
    .C1(_2575_),
    .X(_2576_));
 sky130_fd_sc_hd__a21o_2 _5828_ (.A1(_2504_),
    .A2(_2564_),
    .B1(_2576_),
    .X(alu_out[7]));
 sky130_fd_sc_hd__inv_2 _5829_ (.A(_2418_),
    .Y(_2577_));
 sky130_fd_sc_hd__mux2_2 _5830_ (.A0(_2577_),
    .A1(_2498_),
    .S(_1803_),
    .X(_2578_));
 sky130_fd_sc_hd__inv_2 _5831_ (.A(_2578_),
    .Y(_2579_));
 sky130_fd_sc_hd__inv_2 _5832_ (.A(_2287_),
    .Y(_2580_));
 sky130_fd_sc_hd__mux2_2 _5833_ (.A0(_2230_),
    .A1(_2580_),
    .S(_1839_),
    .X(_2581_));
 sky130_fd_sc_hd__inv_2 _5834_ (.A(_2581_),
    .Y(_2582_));
 sky130_fd_sc_hd__mux2_2 _5835_ (.A0(_2547_),
    .A1(_2582_),
    .S(_2363_),
    .X(_2583_));
 sky130_fd_sc_hd__mux2_2 _5836_ (.A0(_2579_),
    .A1(_2583_),
    .S(_2252_),
    .X(_2584_));
 sky130_fd_sc_hd__or3b_2 _5837_ (.A(_1758_),
    .B(_2331_),
    .C_N(_1148_),
    .X(_2585_));
 sky130_fd_sc_hd__o2bb2a_2 _5838_ (.A1_N(_2105_),
    .A2_N(_2584_),
    .B1(_2487_),
    .B2(_2585_),
    .X(_2586_));
 sky130_fd_sc_hd__nor2_2 _5839_ (.A(_2335_),
    .B(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__nand2_2 _5840_ (.A(_2040_),
    .B(_2372_),
    .Y(_2588_));
 sky130_fd_sc_hd__o21ai_2 _5841_ (.A1(_1880_),
    .A2(_2588_),
    .B1(_2421_),
    .Y(_2589_));
 sky130_fd_sc_hd__or2_2 _5842_ (.A(_1666_),
    .B(_2040_),
    .X(_2590_));
 sky130_fd_sc_hd__nor2_2 _5843_ (.A(_2039_),
    .B(_2102_),
    .Y(_2591_));
 sky130_fd_sc_hd__a2bb2o_2 _5844_ (.A1_N(_2038_),
    .A2_N(_2590_),
    .B1(_2591_),
    .B2(_2253_),
    .X(_2592_));
 sky130_fd_sc_hd__nand4_2 _5845_ (.A(_1111_),
    .B(_1125_),
    .C(_1145_),
    .D(_1166_),
    .Y(_2593_));
 sky130_fd_sc_hd__nand2_2 _5846_ (.A(_1060_),
    .B(_1083_),
    .Y(_2594_));
 sky130_fd_sc_hd__nand2_2 _5847_ (.A(opcode[0]),
    .B(_2503_),
    .Y(_2595_));
 sky130_fd_sc_hd__o31a_2 _5848_ (.A1(_1416_),
    .A2(_2593_),
    .A3(_2594_),
    .B1(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__xor2_2 _5849_ (.A(_1528_),
    .B(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__xor2_2 _5850_ (.A(_2229_),
    .B(_2597_),
    .X(_2598_));
 sky130_fd_sc_hd__a21oi_2 _5851_ (.A1(_2562_),
    .A2(_2560_),
    .B1(_2559_),
    .Y(_2599_));
 sky130_fd_sc_hd__a311o_2 _5852_ (.A1(_2511_),
    .A2(_2512_),
    .A3(_2518_),
    .B1(_2542_),
    .C1(_2599_),
    .X(_2600_));
 sky130_fd_sc_hd__o21ai_2 _5853_ (.A1(_2539_),
    .A2(_2559_),
    .B1(_2560_),
    .Y(_2601_));
 sky130_fd_sc_hd__nand2_2 _5854_ (.A(_2600_),
    .B(_2601_),
    .Y(_2602_));
 sky130_fd_sc_hd__xnor2_2 _5855_ (.A(_2598_),
    .B(_2602_),
    .Y(_2603_));
 sky130_fd_sc_hd__o32a_2 _5856_ (.A1(_2587_),
    .A2(_2589_),
    .A3(_2592_),
    .B1(_2603_),
    .B2(_2408_),
    .X(alu_out[8]));
 sky130_fd_sc_hd__nor2_2 _5857_ (.A(_2390_),
    .B(_2590_),
    .Y(_2604_));
 sky130_fd_sc_hd__nor2_2 _5858_ (.A(_1111_),
    .B(_2102_),
    .Y(_2605_));
 sky130_fd_sc_hd__a22o_2 _5859_ (.A1(_2404_),
    .A2(_2605_),
    .B1(_2591_),
    .B2(_2356_),
    .X(_2606_));
 sky130_fd_sc_hd__or3_2 _5860_ (.A(_2504_),
    .B(_2604_),
    .C(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__mux2_2 _5861_ (.A0(_2457_),
    .A1(_2525_),
    .S(_1877_),
    .X(_2608_));
 sky130_fd_sc_hd__and2_2 _5862_ (.A(_2353_),
    .B(_2358_),
    .X(_2609_));
 sky130_fd_sc_hd__mux2_2 _5863_ (.A0(_2565_),
    .A1(_2609_),
    .S(_1803_),
    .X(_2610_));
 sky130_fd_sc_hd__nand2_2 _5864_ (.A(_2252_),
    .B(_2610_),
    .Y(_2611_));
 sky130_fd_sc_hd__o21ai_2 _5865_ (.A1(_2426_),
    .A2(_2608_),
    .B1(_2611_),
    .Y(_2612_));
 sky130_fd_sc_hd__a2bb2o_2 _5866_ (.A1_N(_2340_),
    .A2_N(_2487_),
    .B1(_2612_),
    .B2(_2530_),
    .X(_2613_));
 sky130_fd_sc_hd__and2_2 _5867_ (.A(_1087_),
    .B(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__o41a_2 _5868_ (.A1(_1528_),
    .A2(_1416_),
    .A3(_2593_),
    .A4(_2594_),
    .B1(_2595_),
    .X(_2615_));
 sky130_fd_sc_hd__xnor2_2 _5869_ (.A(_1542_),
    .B(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__xor2_2 _5870_ (.A(_2246_),
    .B(_2616_),
    .X(_2617_));
 sky130_fd_sc_hd__and2_2 _5871_ (.A(_2600_),
    .B(_2601_),
    .X(_2618_));
 sky130_fd_sc_hd__a2bb2o_2 _5872_ (.A1_N(_2229_),
    .A2_N(_2597_),
    .B1(_2598_),
    .B2(_2618_),
    .X(_2619_));
 sky130_fd_sc_hd__xor2_2 _5873_ (.A(_2617_),
    .B(_2619_),
    .X(_2620_));
 sky130_fd_sc_hd__buf_1 _5874_ (.A(_2333_),
    .X(_2621_));
 sky130_fd_sc_hd__o22a_2 _5875_ (.A1(_2607_),
    .A2(_2614_),
    .B1(_2620_),
    .B2(_2621_),
    .X(alu_out[9]));
 sky130_fd_sc_hd__o21a_2 _5876_ (.A1(_1839_),
    .A2(_2211_),
    .B1(_2248_),
    .X(_2622_));
 sky130_fd_sc_hd__mux2_2 _5877_ (.A0(_2581_),
    .A1(_2622_),
    .S(_1146_),
    .X(_2623_));
 sky130_fd_sc_hd__inv_2 _5878_ (.A(_2623_),
    .Y(_2624_));
 sky130_fd_sc_hd__mux2_2 _5879_ (.A0(_2548_),
    .A1(_2624_),
    .S(_2426_),
    .X(_2625_));
 sky130_fd_sc_hd__a22oi_2 _5880_ (.A1(_2546_),
    .A2(_2570_),
    .B1(_2625_),
    .B2(_2105_),
    .Y(_2626_));
 sky130_fd_sc_hd__nor2_2 _5881_ (.A(_2335_),
    .B(_2626_),
    .Y(_2627_));
 sky130_fd_sc_hd__o22ai_2 _5882_ (.A1(_2441_),
    .A2(_2588_),
    .B1(_2590_),
    .B2(_2444_),
    .Y(_2628_));
 sky130_fd_sc_hd__a211o_2 _5883_ (.A1(_2427_),
    .A2(_2591_),
    .B1(_2628_),
    .C1(_2504_),
    .X(_2629_));
 sky130_fd_sc_hd__or2b_2 _5884_ (.A(_1528_),
    .B_N(_1542_),
    .X(_2630_));
 sky130_fd_sc_hd__o41a_2 _5885_ (.A1(_2630_),
    .A2(_1416_),
    .A3(_2593_),
    .A4(_2594_),
    .B1(_2595_),
    .X(_2631_));
 sky130_fd_sc_hd__xnor2_2 _5886_ (.A(_1558_),
    .B(_2631_),
    .Y(_2632_));
 sky130_fd_sc_hd__xor2_2 _5887_ (.A(_2210_),
    .B(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__o22a_2 _5888_ (.A1(_2229_),
    .A2(_2597_),
    .B1(_2616_),
    .B2(_2246_),
    .X(_2634_));
 sky130_fd_sc_hd__a21oi_2 _5889_ (.A1(_2246_),
    .A2(_2616_),
    .B1(_2634_),
    .Y(_2635_));
 sky130_fd_sc_hd__a31o_2 _5890_ (.A1(_2598_),
    .A2(_2618_),
    .A3(_2617_),
    .B1(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__xor2_2 _5891_ (.A(_2633_),
    .B(_2636_),
    .X(_2637_));
 sky130_fd_sc_hd__o22a_2 _5892_ (.A1(_2627_),
    .A2(_2629_),
    .B1(_2637_),
    .B2(_2621_),
    .X(alu_out[10]));
 sky130_fd_sc_hd__nand3b_2 _5893_ (.A_N(_1528_),
    .B(_1542_),
    .C(_1558_),
    .Y(_2638_));
 sky130_fd_sc_hd__or4_2 _5894_ (.A(_2638_),
    .B(_1416_),
    .C(_2593_),
    .D(_2594_),
    .X(_2639_));
 sky130_fd_sc_hd__nand3_2 _5895_ (.A(_1572_),
    .B(_2595_),
    .C(_2639_),
    .Y(_2640_));
 sky130_fd_sc_hd__a21o_2 _5896_ (.A1(_2595_),
    .A2(_2639_),
    .B1(_1572_),
    .X(_2641_));
 sky130_fd_sc_hd__a21o_2 _5897_ (.A1(_2640_),
    .A2(_2641_),
    .B1(_2193_),
    .X(_2642_));
 sky130_fd_sc_hd__nand3_2 _5898_ (.A(_2193_),
    .B(_2640_),
    .C(_2641_),
    .Y(_2643_));
 sky130_fd_sc_hd__nand2_2 _5899_ (.A(_2642_),
    .B(_2643_),
    .Y(_2644_));
 sky130_fd_sc_hd__nor2_2 _5900_ (.A(_2210_),
    .B(_2632_),
    .Y(_2645_));
 sky130_fd_sc_hd__a21oi_2 _5901_ (.A1(_2633_),
    .A2(_2636_),
    .B1(_2645_),
    .Y(_2646_));
 sky130_fd_sc_hd__xnor2_2 _5902_ (.A(_2644_),
    .B(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__inv_2 _5903_ (.A(_2567_),
    .Y(_2648_));
 sky130_fd_sc_hd__and2_2 _5904_ (.A(_2352_),
    .B(_2350_),
    .X(_2649_));
 sky130_fd_sc_hd__mux2_2 _5905_ (.A0(_2609_),
    .A1(_2649_),
    .S(_1803_),
    .X(_2650_));
 sky130_fd_sc_hd__mux2_2 _5906_ (.A0(_2648_),
    .A1(_2650_),
    .S(_2501_),
    .X(_2651_));
 sky130_fd_sc_hd__a2bb2o_2 _5907_ (.A1_N(_2458_),
    .A2_N(_2487_),
    .B1(_2651_),
    .B2(_2530_),
    .X(_2652_));
 sky130_fd_sc_hd__and2_2 _5908_ (.A(_1087_),
    .B(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__a31o_2 _5909_ (.A1(_2468_),
    .A2(_2530_),
    .A3(_2475_),
    .B1(_2503_),
    .X(_2654_));
 sky130_fd_sc_hd__a22o_2 _5910_ (.A1(_2471_),
    .A2(_2605_),
    .B1(_2591_),
    .B2(_2462_),
    .X(_2655_));
 sky130_fd_sc_hd__or2_2 _5911_ (.A(_2654_),
    .B(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__o2bb2a_2 _5912_ (.A1_N(_2504_),
    .A2_N(_2647_),
    .B1(_2653_),
    .B2(_2656_),
    .X(alu_out[11]));
 sky130_fd_sc_hd__and4b_2 _5913_ (.A_N(_1416_),
    .B(_1573_),
    .C(_2506_),
    .D(_2535_),
    .X(_2657_));
 sky130_fd_sc_hd__buf_1 _5914_ (.A(_2657_),
    .X(_2658_));
 sky130_fd_sc_hd__or3_2 _5915_ (.A(_1464_),
    .B(_2536_),
    .C(_2658_),
    .X(_2659_));
 sky130_fd_sc_hd__o21ai_2 _5916_ (.A1(_2536_),
    .A2(_2658_),
    .B1(_1464_),
    .Y(_2660_));
 sky130_fd_sc_hd__a21o_2 _5917_ (.A1(_2659_),
    .A2(_2660_),
    .B1(_2175_),
    .X(_2661_));
 sky130_fd_sc_hd__nand3_2 _5918_ (.A(_2175_),
    .B(_2659_),
    .C(_2660_),
    .Y(_2662_));
 sky130_fd_sc_hd__nand2_2 _5919_ (.A(_2661_),
    .B(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__and3_2 _5920_ (.A(_2633_),
    .B(_2642_),
    .C(_2643_),
    .X(_2664_));
 sky130_fd_sc_hd__nand3_2 _5921_ (.A(_2598_),
    .B(_2617_),
    .C(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__and3_2 _5922_ (.A(_2193_),
    .B(_2640_),
    .C(_2641_),
    .X(_2666_));
 sky130_fd_sc_hd__a221oi_2 _5923_ (.A1(_2645_),
    .A2(_2642_),
    .B1(_2664_),
    .B2(_2635_),
    .C1(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__o21a_2 _5924_ (.A1(_2602_),
    .A2(_2665_),
    .B1(_2667_),
    .X(_2668_));
 sky130_fd_sc_hd__or2_2 _5925_ (.A(_2663_),
    .B(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__nand2_2 _5926_ (.A(_2663_),
    .B(_2668_),
    .Y(_2670_));
 sky130_fd_sc_hd__nand2_2 _5927_ (.A(_2669_),
    .B(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__nor2_2 _5928_ (.A(_2428_),
    .B(_2288_),
    .Y(_2672_));
 sky130_fd_sc_hd__mux2_2 _5929_ (.A0(_2547_),
    .A1(_2672_),
    .S(_1147_),
    .X(_2673_));
 sky130_fd_sc_hd__nor2_2 _5930_ (.A(_2212_),
    .B(_2429_),
    .Y(_2674_));
 sky130_fd_sc_hd__o21a_2 _5931_ (.A1(_1800_),
    .A2(_2194_),
    .B1(_2176_),
    .X(_2675_));
 sky130_fd_sc_hd__mux2_2 _5932_ (.A0(_2674_),
    .A1(_2675_),
    .S(_1147_),
    .X(_2676_));
 sky130_fd_sc_hd__mux2_2 _5933_ (.A0(_2673_),
    .A1(_2676_),
    .S(_2501_),
    .X(_2677_));
 sky130_fd_sc_hd__mux2_2 _5934_ (.A0(_2502_),
    .A1(_2677_),
    .S(_2104_),
    .X(_2678_));
 sky130_fd_sc_hd__or3b_2 _5935_ (.A(_1666_),
    .B(_2039_),
    .C_N(_2251_),
    .X(_2679_));
 sky130_fd_sc_hd__o221a_2 _5936_ (.A1(_2486_),
    .A2(_2588_),
    .B1(_2679_),
    .B2(_1962_),
    .C1(_2333_),
    .X(_2680_));
 sky130_fd_sc_hd__a21bo_2 _5937_ (.A1(_2491_),
    .A2(_2591_),
    .B1_N(_2680_),
    .X(_2681_));
 sky130_fd_sc_hd__a21oi_2 _5938_ (.A1(_1087_),
    .A2(_2678_),
    .B1(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__a21oi_2 _5939_ (.A1(_2504_),
    .A2(_2671_),
    .B1(_2682_),
    .Y(alu_out[12]));
 sky130_fd_sc_hd__inv_2 _5940_ (.A(_1480_),
    .Y(_2683_));
 sky130_fd_sc_hd__a211o_2 _5941_ (.A1(_1464_),
    .A2(_2657_),
    .B1(_2411_),
    .C1(_2683_),
    .X(_2684_));
 sky130_fd_sc_hd__or2_2 _5942_ (.A(_1464_),
    .B(_2411_),
    .X(_2685_));
 sky130_fd_sc_hd__o211ai_2 _5943_ (.A1(_2536_),
    .A2(_2657_),
    .B1(_2685_),
    .C1(_2683_),
    .Y(_2686_));
 sky130_fd_sc_hd__and3_2 _5944_ (.A(_2160_),
    .B(_2684_),
    .C(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__a21oi_2 _5945_ (.A1(_2684_),
    .A2(_2686_),
    .B1(_2160_),
    .Y(_2688_));
 sky130_fd_sc_hd__or2_2 _5946_ (.A(_2687_),
    .B(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__and3b_2 _5947_ (.A_N(_2689_),
    .B(_2669_),
    .C(_2661_),
    .X(_2690_));
 sky130_fd_sc_hd__a21boi_2 _5948_ (.A1(_2661_),
    .A2(_2669_),
    .B1_N(_2689_),
    .Y(_2691_));
 sky130_fd_sc_hd__mux2_2 _5949_ (.A0(_2378_),
    .A1(_2381_),
    .S(_2178_),
    .X(_2692_));
 sky130_fd_sc_hd__nor2_2 _5950_ (.A(_2692_),
    .B(_2679_),
    .Y(_2693_));
 sky130_fd_sc_hd__a22o_2 _5951_ (.A1(_2522_),
    .A2(_2605_),
    .B1(_2591_),
    .B2(_2531_),
    .X(_2694_));
 sky130_fd_sc_hd__or3_2 _5952_ (.A(_2503_),
    .B(_2693_),
    .C(_2694_),
    .X(_2695_));
 sky130_fd_sc_hd__mux2_2 _5953_ (.A0(_2340_),
    .A1(_2608_),
    .S(_1879_),
    .X(_2696_));
 sky130_fd_sc_hd__and2_2 _5954_ (.A(_2345_),
    .B(_2349_),
    .X(_2697_));
 sky130_fd_sc_hd__mux2_2 _5955_ (.A0(_2649_),
    .A1(_2697_),
    .S(_1803_),
    .X(_2698_));
 sky130_fd_sc_hd__mux2_2 _5956_ (.A0(_2610_),
    .A1(_2698_),
    .S(_2251_),
    .X(_2699_));
 sky130_fd_sc_hd__nand2_2 _5957_ (.A(_2104_),
    .B(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__o21a_2 _5958_ (.A1(_2104_),
    .A2(_2696_),
    .B1(_2700_),
    .X(_2701_));
 sky130_fd_sc_hd__nor2_2 _5959_ (.A(_2335_),
    .B(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__o32a_2 _5960_ (.A1(_2421_),
    .A2(_2690_),
    .A3(_2691_),
    .B1(_2695_),
    .B2(_2702_),
    .X(alu_out[13]));
 sky130_fd_sc_hd__nor2_2 _5961_ (.A(_2161_),
    .B(_2142_),
    .Y(_2703_));
 sky130_fd_sc_hd__mux2_2 _5962_ (.A0(_2675_),
    .A1(_2703_),
    .S(_2347_),
    .X(_2704_));
 sky130_fd_sc_hd__mux2_2 _5963_ (.A0(_2624_),
    .A1(_2704_),
    .S(_2501_),
    .X(_2705_));
 sky130_fd_sc_hd__mux2_2 _5964_ (.A0(_2549_),
    .A1(_2705_),
    .S(_2104_),
    .X(_2706_));
 sky130_fd_sc_hd__and2_2 _5965_ (.A(_1087_),
    .B(_2706_),
    .X(_2707_));
 sky130_fd_sc_hd__o221a_2 _5966_ (.A1(_2553_),
    .A2(_2588_),
    .B1(_2679_),
    .B2(_2442_),
    .C1(_2333_),
    .X(_2708_));
 sky130_fd_sc_hd__a21bo_2 _5967_ (.A1(_2550_),
    .A2(_2591_),
    .B1_N(_2708_),
    .X(_2709_));
 sky130_fd_sc_hd__a31o_2 _5968_ (.A1(_1464_),
    .A2(_1480_),
    .A3(_2657_),
    .B1(_2411_),
    .X(_2710_));
 sky130_fd_sc_hd__xor2_2 _5969_ (.A(_1494_),
    .B(_2710_),
    .X(_2711_));
 sky130_fd_sc_hd__xnor2_2 _5970_ (.A(_2140_),
    .B(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__o21ba_2 _5971_ (.A1(_2661_),
    .A2(_2688_),
    .B1_N(_2687_),
    .X(_2713_));
 sky130_fd_sc_hd__o21ai_2 _5972_ (.A1(_2669_),
    .A2(_2689_),
    .B1(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__xnor2_2 _5973_ (.A(_2712_),
    .B(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__o22a_2 _5974_ (.A1(_2707_),
    .A2(_2709_),
    .B1(_2715_),
    .B2(_2621_),
    .X(alu_out[14]));
 sky130_fd_sc_hd__and2_2 _5975_ (.A(_2573_),
    .B(_2591_),
    .X(_2716_));
 sky130_fd_sc_hd__and2_2 _5976_ (.A(_2344_),
    .B(_2342_),
    .X(_2717_));
 sky130_fd_sc_hd__mux2_2 _5977_ (.A0(_2697_),
    .A1(_2717_),
    .S(_1803_),
    .X(_2718_));
 sky130_fd_sc_hd__mux2_2 _5978_ (.A0(_2650_),
    .A1(_2718_),
    .S(_2251_),
    .X(_2719_));
 sky130_fd_sc_hd__mux2_2 _5979_ (.A0(_2569_),
    .A1(_2719_),
    .S(_2104_),
    .X(_2720_));
 sky130_fd_sc_hd__a41o_2 _5980_ (.A1(_2468_),
    .A2(_2530_),
    .A3(_2426_),
    .A4(_2472_),
    .B1(_2503_),
    .X(_2721_));
 sky130_fd_sc_hd__a221o_2 _5981_ (.A1(_2571_),
    .A2(_2605_),
    .B1(_2720_),
    .B2(_1087_),
    .C1(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__a21oi_2 _5982_ (.A1(_1495_),
    .A2(_2657_),
    .B1(_2536_),
    .Y(_2723_));
 sky130_fd_sc_hd__xnor2_2 _5983_ (.A(_1511_),
    .B(_2723_),
    .Y(_2724_));
 sky130_fd_sc_hd__xnor2_2 _5984_ (.A(_2123_),
    .B(_2724_),
    .Y(_2725_));
 sky130_fd_sc_hd__or2_2 _5985_ (.A(_2140_),
    .B(_2711_),
    .X(_2726_));
 sky130_fd_sc_hd__or2b_2 _5986_ (.A(_2712_),
    .B_N(_2714_),
    .X(_2727_));
 sky130_fd_sc_hd__nand2_2 _5987_ (.A(_2726_),
    .B(_2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__xnor2_2 _5988_ (.A(_2725_),
    .B(_2728_),
    .Y(_2729_));
 sky130_fd_sc_hd__o22a_2 _5989_ (.A1(_2716_),
    .A2(_2722_),
    .B1(_2729_),
    .B2(_2621_),
    .X(alu_out[15]));
 sky130_fd_sc_hd__nor2_2 _5990_ (.A(_2041_),
    .B(_2102_),
    .Y(_2730_));
 sky130_fd_sc_hd__nor2_2 _5991_ (.A(_1111_),
    .B(_2335_),
    .Y(_2731_));
 sky130_fd_sc_hd__nor2_2 _5992_ (.A(_2347_),
    .B(_2622_),
    .Y(_2732_));
 sky130_fd_sc_hd__a21o_2 _5993_ (.A1(_2327_),
    .A2(_2675_),
    .B1(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__o21a_2 _5994_ (.A1(_1169_),
    .A2(_2124_),
    .B1(_1875_),
    .X(_2734_));
 sky130_fd_sc_hd__mux2_2 _5995_ (.A0(_2703_),
    .A1(_2734_),
    .S(_2347_),
    .X(_2735_));
 sky130_fd_sc_hd__mux2_2 _5996_ (.A0(_2733_),
    .A1(_2735_),
    .S(_1879_),
    .X(_2736_));
 sky130_fd_sc_hd__nor2b_2 _5997_ (.A(_1060_),
    .B_N(_1085_),
    .Y(_2737_));
 sky130_fd_sc_hd__nand2_2 _5998_ (.A(_1127_),
    .B(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__o21ai_2 _5999_ (.A1(_2585_),
    .A2(_2738_),
    .B1(_2333_),
    .Y(_2739_));
 sky130_fd_sc_hd__a221o_2 _6000_ (.A1(_2584_),
    .A2(_2731_),
    .B1(_2736_),
    .B2(_2496_),
    .C1(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__buf_1 _6001_ (.A(_2536_),
    .X(_2741_));
 sky130_fd_sc_hd__a21oi_2 _6002_ (.A1(_1512_),
    .A2(_2658_),
    .B1(_2741_),
    .Y(_2742_));
 sky130_fd_sc_hd__xnor2_2 _6003_ (.A(_1587_),
    .B(_2742_),
    .Y(_2743_));
 sky130_fd_sc_hd__xor2_2 _6004_ (.A(_1874_),
    .B(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__or4_2 _6005_ (.A(_2663_),
    .B(_2689_),
    .C(_2712_),
    .D(_2725_),
    .X(_2745_));
 sky130_fd_sc_hd__or3_2 _6006_ (.A(_2712_),
    .B(_2713_),
    .C(_2725_),
    .X(_2746_));
 sky130_fd_sc_hd__a21o_2 _6007_ (.A1(_2123_),
    .A2(_2724_),
    .B1(_2726_),
    .X(_2747_));
 sky130_fd_sc_hd__o211a_2 _6008_ (.A1(_2123_),
    .A2(_2724_),
    .B1(_2746_),
    .C1(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__o21ai_2 _6009_ (.A1(_2668_),
    .A2(_2745_),
    .B1(_2748_),
    .Y(_2749_));
 sky130_fd_sc_hd__xor2_2 _6010_ (.A(_2744_),
    .B(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__o22a_2 _6011_ (.A1(_2730_),
    .A2(_2740_),
    .B1(_2750_),
    .B2(_2621_),
    .X(alu_out[16]));
 sky130_fd_sc_hd__mux2_2 _6012_ (.A0(_2649_),
    .A1(_2697_),
    .S(_2327_),
    .X(_2751_));
 sky130_fd_sc_hd__nor2_2 _6013_ (.A(_2341_),
    .B(_2401_),
    .Y(_2752_));
 sky130_fd_sc_hd__mux2_2 _6014_ (.A0(_2717_),
    .A1(_2752_),
    .S(_1146_),
    .X(_2753_));
 sky130_fd_sc_hd__mux2_2 _6015_ (.A0(_2751_),
    .A1(_2753_),
    .S(_2252_),
    .X(_2754_));
 sky130_fd_sc_hd__and2_2 _6016_ (.A(_2496_),
    .B(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__mux2_2 _6017_ (.A0(_2565_),
    .A1(_2609_),
    .S(_1148_),
    .X(_2756_));
 sky130_fd_sc_hd__mux2_2 _6018_ (.A0(_2527_),
    .A1(_2756_),
    .S(_2426_),
    .X(_2757_));
 sky130_fd_sc_hd__a31o_2 _6019_ (.A1(_1127_),
    .A2(_2524_),
    .A3(_2737_),
    .B1(_2503_),
    .X(_2758_));
 sky130_fd_sc_hd__nor2_2 _6020_ (.A(_2102_),
    .B(_2406_),
    .Y(_2759_));
 sky130_fd_sc_hd__a211o_2 _6021_ (.A1(_2757_),
    .A2(_2731_),
    .B1(_2758_),
    .C1(_2759_),
    .X(_2760_));
 sky130_fd_sc_hd__a31o_2 _6022_ (.A1(_1512_),
    .A2(_1587_),
    .A3(_2658_),
    .B1(_2741_),
    .X(_2761_));
 sky130_fd_sc_hd__xor2_2 _6023_ (.A(_1601_),
    .B(_2761_),
    .X(_2762_));
 sky130_fd_sc_hd__xor2_2 _6024_ (.A(_1858_),
    .B(_2762_),
    .X(_2763_));
 sky130_fd_sc_hd__nor2_2 _6025_ (.A(_1874_),
    .B(_2743_),
    .Y(_2764_));
 sky130_fd_sc_hd__a21oi_2 _6026_ (.A1(_2744_),
    .A2(_2749_),
    .B1(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__xnor2_2 _6027_ (.A(_2763_),
    .B(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__o22a_2 _6028_ (.A1(_2755_),
    .A2(_2760_),
    .B1(_2766_),
    .B2(_2621_),
    .X(alu_out[17]));
 sky130_fd_sc_hd__a31o_2 _6029_ (.A1(_1512_),
    .A2(_1602_),
    .A3(_2658_),
    .B1(_2536_),
    .X(_2767_));
 sky130_fd_sc_hd__xor2_2 _6030_ (.A(_1634_),
    .B(_2767_),
    .X(_2768_));
 sky130_fd_sc_hd__xnor2_2 _6031_ (.A(_1820_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__nand2_2 _6032_ (.A(_2744_),
    .B(_2763_),
    .Y(_2770_));
 sky130_fd_sc_hd__inv_2 _6033_ (.A(_2770_),
    .Y(_2771_));
 sky130_fd_sc_hd__o22a_2 _6034_ (.A1(_1874_),
    .A2(_2743_),
    .B1(_2762_),
    .B2(_1858_),
    .X(_2772_));
 sky130_fd_sc_hd__a21o_2 _6035_ (.A1(_1858_),
    .A2(_2762_),
    .B1(_2772_),
    .X(_2773_));
 sky130_fd_sc_hd__a21bo_2 _6036_ (.A1(_2749_),
    .A2(_2771_),
    .B1_N(_2773_),
    .X(_2774_));
 sky130_fd_sc_hd__xnor2_2 _6037_ (.A(_2769_),
    .B(_2774_),
    .Y(_2775_));
 sky130_fd_sc_hd__nor2_2 _6038_ (.A(_2102_),
    .B(_2445_),
    .Y(_2776_));
 sky130_fd_sc_hd__o21a_2 _6039_ (.A1(_1669_),
    .A2(_1821_),
    .B1(_1860_),
    .X(_2777_));
 sky130_fd_sc_hd__mux2_2 _6040_ (.A0(_2734_),
    .A1(_2777_),
    .S(_1877_),
    .X(_2778_));
 sky130_fd_sc_hd__mux2_2 _6041_ (.A0(_2704_),
    .A1(_2778_),
    .S(_1879_),
    .X(_2779_));
 sky130_fd_sc_hd__o21ai_2 _6042_ (.A1(_2420_),
    .A2(_2738_),
    .B1(_2333_),
    .Y(_2780_));
 sky130_fd_sc_hd__a221o_2 _6043_ (.A1(_2625_),
    .A2(_2731_),
    .B1(_2779_),
    .B2(_2496_),
    .C1(_2780_),
    .X(_2781_));
 sky130_fd_sc_hd__o22a_2 _6044_ (.A1(_2408_),
    .A2(_2775_),
    .B1(_2776_),
    .B2(_2781_),
    .X(alu_out[18]));
 sky130_fd_sc_hd__a41o_2 _6045_ (.A1(_1512_),
    .A2(_1602_),
    .A3(_1634_),
    .A4(_2658_),
    .B1(_2536_),
    .X(_2782_));
 sky130_fd_sc_hd__xor2_2 _6046_ (.A(_1618_),
    .B(_2782_),
    .X(_2783_));
 sky130_fd_sc_hd__xnor2_2 _6047_ (.A(_1838_),
    .B(_2783_),
    .Y(_2784_));
 sky130_fd_sc_hd__nand2_2 _6048_ (.A(_1820_),
    .B(_2768_),
    .Y(_2785_));
 sky130_fd_sc_hd__nor2_2 _6049_ (.A(_1820_),
    .B(_2768_),
    .Y(_2786_));
 sky130_fd_sc_hd__a21oi_2 _6050_ (.A1(_2785_),
    .A2(_2774_),
    .B1(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__xnor2_2 _6051_ (.A(_2784_),
    .B(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__nor2_2 _6052_ (.A(_2421_),
    .B(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__o21a_2 _6053_ (.A1(_1800_),
    .A2(_1821_),
    .B1(_2399_),
    .X(_2790_));
 sky130_fd_sc_hd__mux2_2 _6054_ (.A0(_2752_),
    .A1(_2790_),
    .S(_1147_),
    .X(_2791_));
 sky130_fd_sc_hd__mux2_2 _6055_ (.A0(_2718_),
    .A1(_2791_),
    .S(_2501_),
    .X(_2792_));
 sky130_fd_sc_hd__nor2_2 _6056_ (.A(_2458_),
    .B(_2738_),
    .Y(_2793_));
 sky130_fd_sc_hd__a221o_2 _6057_ (.A1(_2651_),
    .A2(_2731_),
    .B1(_2792_),
    .B2(_2496_),
    .C1(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__a211o_2 _6058_ (.A1(_2373_),
    .A2(_2476_),
    .B1(_2789_),
    .C1(_2794_),
    .X(alu_out[19]));
 sky130_fd_sc_hd__nor2_2 _6059_ (.A(_2102_),
    .B(_2488_),
    .Y(_2795_));
 sky130_fd_sc_hd__mux2_2 _6060_ (.A0(_2585_),
    .A1(_2578_),
    .S(_2426_),
    .X(_2796_));
 sky130_fd_sc_hd__inv_2 _6061_ (.A(_2737_),
    .Y(_2797_));
 sky130_fd_sc_hd__o31ai_2 _6062_ (.A1(_2040_),
    .A2(_2796_),
    .A3(_2797_),
    .B1(_2421_),
    .Y(_2798_));
 sky130_fd_sc_hd__mux2_2 _6063_ (.A0(_2583_),
    .A1(_2733_),
    .S(_2426_),
    .X(_2799_));
 sky130_fd_sc_hd__and2b_2 _6064_ (.A_N(_1840_),
    .B(_1801_),
    .X(_2800_));
 sky130_fd_sc_hd__mux2_2 _6065_ (.A0(_2777_),
    .A1(_2800_),
    .S(_1147_),
    .X(_2801_));
 sky130_fd_sc_hd__mux2_2 _6066_ (.A0(_2735_),
    .A1(_2801_),
    .S(_2252_),
    .X(_2802_));
 sky130_fd_sc_hd__a22o_2 _6067_ (.A1(_2799_),
    .A2(_2731_),
    .B1(_2802_),
    .B2(_2496_),
    .X(_2803_));
 sky130_fd_sc_hd__a31o_2 _6068_ (.A1(_1512_),
    .A2(_1635_),
    .A3(_2658_),
    .B1(_2536_),
    .X(_2804_));
 sky130_fd_sc_hd__xor2_2 _6069_ (.A(_1256_),
    .B(_2804_),
    .X(_2805_));
 sky130_fd_sc_hd__nor2_2 _6070_ (.A(_1798_),
    .B(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__and2_2 _6071_ (.A(_1798_),
    .B(_2805_),
    .X(_2807_));
 sky130_fd_sc_hd__or2_2 _6072_ (.A(_2806_),
    .B(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__or2_2 _6073_ (.A(_2769_),
    .B(_2784_),
    .X(_2809_));
 sky130_fd_sc_hd__a211o_2 _6074_ (.A1(_1838_),
    .A2(_2783_),
    .B1(_2768_),
    .C1(_1820_),
    .X(_2810_));
 sky130_fd_sc_hd__or2_2 _6075_ (.A(_1838_),
    .B(_2783_),
    .X(_2811_));
 sky130_fd_sc_hd__o211a_2 _6076_ (.A1(_2773_),
    .A2(_2809_),
    .B1(_2810_),
    .C1(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__inv_2 _6077_ (.A(_2601_),
    .Y(_2813_));
 sky130_fd_sc_hd__or4b_2 _6078_ (.A(_2813_),
    .B(_2665_),
    .C(_2745_),
    .D_N(_2600_),
    .X(_2814_));
 sky130_fd_sc_hd__or2_2 _6079_ (.A(_2667_),
    .B(_2745_),
    .X(_2815_));
 sky130_fd_sc_hd__or2_2 _6080_ (.A(_2770_),
    .B(_2809_),
    .X(_2816_));
 sky130_fd_sc_hd__a31o_2 _6081_ (.A1(_2814_),
    .A2(_2815_),
    .A3(_2748_),
    .B1(_2816_),
    .X(_2817_));
 sky130_fd_sc_hd__nand2_2 _6082_ (.A(_2812_),
    .B(_2817_),
    .Y(_2818_));
 sky130_fd_sc_hd__xnor2_2 _6083_ (.A(_2808_),
    .B(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__o32a_2 _6084_ (.A1(_2795_),
    .A2(_2798_),
    .A3(_2803_),
    .B1(_2819_),
    .B2(_2408_),
    .X(alu_out[20]));
 sky130_fd_sc_hd__nor2_2 _6085_ (.A(_2398_),
    .B(_2395_),
    .Y(_2820_));
 sky130_fd_sc_hd__mux2_2 _6086_ (.A0(_2790_),
    .A1(_2820_),
    .S(_1146_),
    .X(_2821_));
 sky130_fd_sc_hd__mux2_2 _6087_ (.A0(_2753_),
    .A1(_2821_),
    .S(_1126_),
    .X(_2822_));
 sky130_fd_sc_hd__nor2_2 _6088_ (.A(_2040_),
    .B(_2797_),
    .Y(_2823_));
 sky130_fd_sc_hd__mux2_2 _6089_ (.A0(_2756_),
    .A1(_2751_),
    .S(_2426_),
    .X(_2824_));
 sky130_fd_sc_hd__nor2_2 _6090_ (.A(_2102_),
    .B(_2523_),
    .Y(_2825_));
 sky130_fd_sc_hd__a221o_2 _6091_ (.A1(_2528_),
    .A2(_2823_),
    .B1(_2731_),
    .B2(_2824_),
    .C1(_2825_),
    .X(_2826_));
 sky130_fd_sc_hd__a21oi_2 _6092_ (.A1(_2812_),
    .A2(_2817_),
    .B1(_2808_),
    .Y(_2827_));
 sky130_fd_sc_hd__a41o_2 _6093_ (.A1(_1512_),
    .A2(_1256_),
    .A3(_1635_),
    .A4(_2658_),
    .B1(_2741_),
    .X(_2828_));
 sky130_fd_sc_hd__xnor2_2 _6094_ (.A(_1277_),
    .B(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__xor2_2 _6095_ (.A(_1779_),
    .B(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__inv_2 _6096_ (.A(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__nor2_2 _6097_ (.A(_2806_),
    .B(_2827_),
    .Y(_2832_));
 sky130_fd_sc_hd__o21a_2 _6098_ (.A1(_2830_),
    .A2(_2832_),
    .B1(_2503_),
    .X(_2833_));
 sky130_fd_sc_hd__o31a_2 _6099_ (.A1(_2806_),
    .A2(_2827_),
    .A3(_2831_),
    .B1(_2833_),
    .X(_2834_));
 sky130_fd_sc_hd__a211o_2 _6100_ (.A1(_2496_),
    .A2(_2822_),
    .B1(_2826_),
    .C1(_2834_),
    .X(alu_out[21]));
 sky130_fd_sc_hd__and2_2 _6101_ (.A(_1256_),
    .B(_1277_),
    .X(_2835_));
 sky130_fd_sc_hd__a41o_2 _6102_ (.A1(_1512_),
    .A2(_2835_),
    .A3(_1635_),
    .A4(_2658_),
    .B1(_2536_),
    .X(_2836_));
 sky130_fd_sc_hd__xnor2_2 _6103_ (.A(_1446_),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__nand2_2 _6104_ (.A(_1754_),
    .B(_2837_),
    .Y(_2838_));
 sky130_fd_sc_hd__or2_2 _6105_ (.A(_1754_),
    .B(_2837_),
    .X(_2839_));
 sky130_fd_sc_hd__nand2_2 _6106_ (.A(_2838_),
    .B(_2839_),
    .Y(_2840_));
 sky130_fd_sc_hd__or2b_2 _6107_ (.A(_2829_),
    .B_N(_1779_),
    .X(_2841_));
 sky130_fd_sc_hd__and2b_2 _6108_ (.A_N(_1779_),
    .B(_2829_),
    .X(_2842_));
 sky130_fd_sc_hd__a21oi_2 _6109_ (.A1(_2806_),
    .A2(_2841_),
    .B1(_2842_),
    .Y(_2843_));
 sky130_fd_sc_hd__a21boi_2 _6110_ (.A1(_2827_),
    .A2(_2831_),
    .B1_N(_2843_),
    .Y(_2844_));
 sky130_fd_sc_hd__xor2_2 _6111_ (.A(_2840_),
    .B(_2844_),
    .X(_2845_));
 sky130_fd_sc_hd__nor2_2 _6112_ (.A(_2102_),
    .B(_2554_),
    .Y(_2846_));
 sky130_fd_sc_hd__and2_2 _6113_ (.A(_1781_),
    .B(_1756_),
    .X(_2847_));
 sky130_fd_sc_hd__mux2_2 _6114_ (.A0(_2800_),
    .A1(_2847_),
    .S(_1877_),
    .X(_2848_));
 sky130_fd_sc_hd__mux2_2 _6115_ (.A0(_2778_),
    .A1(_2848_),
    .S(_1879_),
    .X(_2849_));
 sky130_fd_sc_hd__a21o_2 _6116_ (.A1(_2495_),
    .A2(_2849_),
    .B1(_2503_),
    .X(_2850_));
 sky130_fd_sc_hd__a221o_2 _6117_ (.A1(_2549_),
    .A2(_2823_),
    .B1(_2731_),
    .B2(_2705_),
    .C1(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__o22a_2 _6118_ (.A1(_2408_),
    .A2(_2845_),
    .B1(_2846_),
    .B2(_2851_),
    .X(alu_out[22]));
 sky130_fd_sc_hd__o21ai_2 _6119_ (.A1(_1446_),
    .A2(_2741_),
    .B1(_2836_),
    .Y(_2852_));
 sky130_fd_sc_hd__xnor2_2 _6120_ (.A(_1430_),
    .B(_2852_),
    .Y(_2853_));
 sky130_fd_sc_hd__xnor2_2 _6121_ (.A(_1731_),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__o21ai_2 _6122_ (.A1(_2840_),
    .A2(_2844_),
    .B1(_2838_),
    .Y(_2855_));
 sky130_fd_sc_hd__xnor2_2 _6123_ (.A(_2854_),
    .B(_2855_),
    .Y(_2856_));
 sky130_fd_sc_hd__nor2_2 _6124_ (.A(_2394_),
    .B(_2392_),
    .Y(_2857_));
 sky130_fd_sc_hd__mux2_2 _6125_ (.A0(_2820_),
    .A1(_2857_),
    .S(_1147_),
    .X(_2858_));
 sky130_fd_sc_hd__mux2_2 _6126_ (.A0(_2791_),
    .A1(_2858_),
    .S(_2501_),
    .X(_2859_));
 sky130_fd_sc_hd__and2_2 _6127_ (.A(_2719_),
    .B(_2731_),
    .X(_2860_));
 sky130_fd_sc_hd__a221o_2 _6128_ (.A1(_2373_),
    .A2(_2572_),
    .B1(_2823_),
    .B2(_2569_),
    .C1(_2860_),
    .X(_2861_));
 sky130_fd_sc_hd__a211o_2 _6129_ (.A1(_2496_),
    .A2(_2859_),
    .B1(_2861_),
    .C1(_2504_),
    .X(_2862_));
 sky130_fd_sc_hd__o21a_2 _6130_ (.A1(_2621_),
    .A2(_2856_),
    .B1(_2862_),
    .X(alu_out[23]));
 sky130_fd_sc_hd__nor2_2 _6131_ (.A(_2586_),
    .B(_2797_),
    .Y(_2863_));
 sky130_fd_sc_hd__nand2_2 _6132_ (.A(_2104_),
    .B(_2373_),
    .Y(_2864_));
 sky130_fd_sc_hd__nor2_2 _6133_ (.A(_2038_),
    .B(_2864_),
    .Y(_2865_));
 sky130_fd_sc_hd__a21oi_2 _6134_ (.A1(_1669_),
    .A2(_1732_),
    .B1(_2035_),
    .Y(_2866_));
 sky130_fd_sc_hd__mux2_2 _6135_ (.A0(_2847_),
    .A1(_2866_),
    .S(_1147_),
    .X(_2867_));
 sky130_fd_sc_hd__o22a_2 _6136_ (.A1(_2254_),
    .A2(_2801_),
    .B1(_2867_),
    .B2(_2336_),
    .X(_2868_));
 sky130_fd_sc_hd__o211a_2 _6137_ (.A1(_2104_),
    .A2(_2736_),
    .B1(_2868_),
    .C1(_1086_),
    .X(_2869_));
 sky130_fd_sc_hd__or3_2 _6138_ (.A(_2504_),
    .B(_2865_),
    .C(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__and4_2 _6139_ (.A(_1512_),
    .B(_2835_),
    .C(_1635_),
    .D(_2658_),
    .X(_2871_));
 sky130_fd_sc_hd__nand2_2 _6140_ (.A(_1447_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__and2_2 _6141_ (.A(_2595_),
    .B(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__xnor2_2 _6142_ (.A(_1384_),
    .B(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__nor2_2 _6143_ (.A(_2033_),
    .B(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__and2_2 _6144_ (.A(_2033_),
    .B(_2874_),
    .X(_2876_));
 sky130_fd_sc_hd__or2_2 _6145_ (.A(_2875_),
    .B(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__or4_2 _6146_ (.A(_2808_),
    .B(_2830_),
    .C(_2840_),
    .D(_2854_),
    .X(_2878_));
 sky130_fd_sc_hd__a311o_2 _6147_ (.A1(_2814_),
    .A2(_2815_),
    .A3(_2748_),
    .B1(_2816_),
    .C1(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a21o_2 _6148_ (.A1(_1731_),
    .A2(_2853_),
    .B1(_2838_),
    .X(_2880_));
 sky130_fd_sc_hd__or2_2 _6149_ (.A(_1731_),
    .B(_2853_),
    .X(_2881_));
 sky130_fd_sc_hd__o311a_2 _6150_ (.A1(_2840_),
    .A2(_2843_),
    .A3(_2854_),
    .B1(_2880_),
    .C1(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__o21a_2 _6151_ (.A1(_2812_),
    .A2(_2878_),
    .B1(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__and3_2 _6152_ (.A(_2877_),
    .B(_2879_),
    .C(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__a21oi_2 _6153_ (.A1(_2879_),
    .A2(_2883_),
    .B1(_2877_),
    .Y(_2885_));
 sky130_fd_sc_hd__nor2_2 _6154_ (.A(_2884_),
    .B(_2885_),
    .Y(_2886_));
 sky130_fd_sc_hd__o22a_2 _6155_ (.A1(_2863_),
    .A2(_2870_),
    .B1(_2886_),
    .B2(_2408_),
    .X(alu_out[24]));
 sky130_fd_sc_hd__or2_2 _6156_ (.A(_2875_),
    .B(_2885_),
    .X(_2887_));
 sky130_fd_sc_hd__a31o_2 _6157_ (.A1(_1447_),
    .A2(_1384_),
    .A3(_2871_),
    .B1(_2741_),
    .X(_2888_));
 sky130_fd_sc_hd__xor2_2 _6158_ (.A(_1370_),
    .B(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__nand2_2 _6159_ (.A(_2015_),
    .B(_2889_),
    .Y(_2890_));
 sky130_fd_sc_hd__inv_2 _6160_ (.A(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__nor2_2 _6161_ (.A(_2015_),
    .B(_2889_),
    .Y(_2892_));
 sky130_fd_sc_hd__or2_2 _6162_ (.A(_2891_),
    .B(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__xnor2_2 _6163_ (.A(_2887_),
    .B(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__nor2_2 _6164_ (.A(_2386_),
    .B(_2391_),
    .Y(_2895_));
 sky130_fd_sc_hd__mux2_2 _6165_ (.A0(_2857_),
    .A1(_2895_),
    .S(_2327_),
    .X(_2896_));
 sky130_fd_sc_hd__o22a_2 _6166_ (.A1(_2255_),
    .A2(_2821_),
    .B1(_2896_),
    .B2(_2337_),
    .X(_2897_));
 sky130_fd_sc_hd__o211a_2 _6167_ (.A1(_2105_),
    .A2(_2754_),
    .B1(_2897_),
    .C1(_1087_),
    .X(_2898_));
 sky130_fd_sc_hd__o21ai_2 _6168_ (.A1(_2390_),
    .A2(_2864_),
    .B1(_2333_),
    .Y(_2899_));
 sky130_fd_sc_hd__a211o_2 _6169_ (.A1(_2613_),
    .A2(_2737_),
    .B1(_2898_),
    .C1(_2899_),
    .X(_2900_));
 sky130_fd_sc_hd__o21a_2 _6170_ (.A1(_2621_),
    .A2(_2894_),
    .B1(_2900_),
    .X(alu_out[25]));
 sky130_fd_sc_hd__inv_2 _6171_ (.A(_1385_),
    .Y(_2901_));
 sky130_fd_sc_hd__a31o_2 _6172_ (.A1(_1447_),
    .A2(_2901_),
    .A3(_2871_),
    .B1(_2741_),
    .X(_2902_));
 sky130_fd_sc_hd__xnor2_2 _6173_ (.A(_1298_),
    .B(_2902_),
    .Y(_2903_));
 sky130_fd_sc_hd__xor2_2 _6174_ (.A(_1996_),
    .B(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__a21oi_2 _6175_ (.A1(_2887_),
    .A2(_2890_),
    .B1(_2892_),
    .Y(_2905_));
 sky130_fd_sc_hd__xnor2_2 _6176_ (.A(_2904_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__nor2_2 _6177_ (.A(_2626_),
    .B(_2797_),
    .Y(_2907_));
 sky130_fd_sc_hd__nor2_2 _6178_ (.A(_2444_),
    .B(_2864_),
    .Y(_2908_));
 sky130_fd_sc_hd__nor2_2 _6179_ (.A(_2017_),
    .B(_1998_),
    .Y(_2909_));
 sky130_fd_sc_hd__mux2_2 _6180_ (.A0(_2866_),
    .A1(_2909_),
    .S(_2327_),
    .X(_2910_));
 sky130_fd_sc_hd__o22a_2 _6181_ (.A1(_2254_),
    .A2(_2848_),
    .B1(_2910_),
    .B2(_2336_),
    .X(_2911_));
 sky130_fd_sc_hd__o211a_2 _6182_ (.A1(_2530_),
    .A2(_2779_),
    .B1(_2911_),
    .C1(_1087_),
    .X(_2912_));
 sky130_fd_sc_hd__or3_2 _6183_ (.A(_2504_),
    .B(_2908_),
    .C(_2912_),
    .X(_2913_));
 sky130_fd_sc_hd__o22a_2 _6184_ (.A1(_2408_),
    .A2(_2906_),
    .B1(_2907_),
    .B2(_2913_),
    .X(alu_out[26]));
 sky130_fd_sc_hd__a41o_2 _6185_ (.A1(_1447_),
    .A2(_1299_),
    .A3(_2901_),
    .A4(_2871_),
    .B1(_2741_),
    .X(_2914_));
 sky130_fd_sc_hd__xor2_2 _6186_ (.A(_1315_),
    .B(_2914_),
    .X(_2915_));
 sky130_fd_sc_hd__or2_2 _6187_ (.A(_1978_),
    .B(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__nand2_2 _6188_ (.A(_1978_),
    .B(_2915_),
    .Y(_2917_));
 sky130_fd_sc_hd__and2_2 _6189_ (.A(_2916_),
    .B(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__o311a_2 _6190_ (.A1(_2875_),
    .A2(_2885_),
    .A3(_2892_),
    .B1(_2904_),
    .C1(_2890_),
    .X(_2919_));
 sky130_fd_sc_hd__o21ba_2 _6191_ (.A1(_1996_),
    .A2(_2903_),
    .B1_N(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__xor2_2 _6192_ (.A(_2918_),
    .B(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__or2_2 _6193_ (.A(_2254_),
    .B(_2858_),
    .X(_2922_));
 sky130_fd_sc_hd__nand2_2 _6194_ (.A(_1669_),
    .B(_1997_),
    .Y(_2923_));
 sky130_fd_sc_hd__nand2_2 _6195_ (.A(_2923_),
    .B(_2384_),
    .Y(_2924_));
 sky130_fd_sc_hd__mux2_2 _6196_ (.A0(_2895_),
    .A1(_2924_),
    .S(_2363_),
    .X(_2925_));
 sky130_fd_sc_hd__o21a_2 _6197_ (.A1(_2337_),
    .A2(_2925_),
    .B1(_1086_),
    .X(_2926_));
 sky130_fd_sc_hd__o211a_2 _6198_ (.A1(_2530_),
    .A2(_2792_),
    .B1(_2922_),
    .C1(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__a221o_2 _6199_ (.A1(_2475_),
    .A2(_2591_),
    .B1(_2652_),
    .B2(_2737_),
    .C1(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__o21bai_2 _6200_ (.A1(_2621_),
    .A2(_2921_),
    .B1_N(_2928_),
    .Y(alu_out[27]));
 sky130_fd_sc_hd__or3_2 _6201_ (.A(_1316_),
    .B(_1385_),
    .C(_2872_),
    .X(_2929_));
 sky130_fd_sc_hd__and2_2 _6202_ (.A(_2595_),
    .B(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__xnor2_2 _6203_ (.A(_1237_),
    .B(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__nor2_2 _6204_ (.A(_1958_),
    .B(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__and2_2 _6205_ (.A(_1958_),
    .B(_2931_),
    .X(_2933_));
 sky130_fd_sc_hd__nor2_2 _6206_ (.A(_2932_),
    .B(_2933_),
    .Y(_2934_));
 sky130_fd_sc_hd__nand2_2 _6207_ (.A(_2904_),
    .B(_2918_),
    .Y(_2935_));
 sky130_fd_sc_hd__nor2_2 _6208_ (.A(_2893_),
    .B(_2935_),
    .Y(_2936_));
 sky130_fd_sc_hd__nor2_2 _6209_ (.A(_2875_),
    .B(_2892_),
    .Y(_2937_));
 sky130_fd_sc_hd__or3b_2 _6210_ (.A(_1996_),
    .B(_2903_),
    .C_N(_2917_),
    .X(_2938_));
 sky130_fd_sc_hd__o311a_2 _6211_ (.A1(_2891_),
    .A2(_2937_),
    .A3(_2935_),
    .B1(_2938_),
    .C1(_2916_),
    .X(_2939_));
 sky130_fd_sc_hd__a21bo_2 _6212_ (.A1(_2885_),
    .A2(_2936_),
    .B1_N(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__xor2_2 _6213_ (.A(_2934_),
    .B(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__nand2_2 _6214_ (.A(_2426_),
    .B(_2591_),
    .Y(_2942_));
 sky130_fd_sc_hd__o21ai_2 _6215_ (.A1(_1962_),
    .A2(_2942_),
    .B1(_2421_),
    .Y(_2943_));
 sky130_fd_sc_hd__nor2_2 _6216_ (.A(_1980_),
    .B(_1960_),
    .Y(_2944_));
 sky130_fd_sc_hd__mux2_2 _6217_ (.A0(_2909_),
    .A1(_2944_),
    .S(_2178_),
    .X(_2945_));
 sky130_fd_sc_hd__o22a_2 _6218_ (.A1(_2255_),
    .A2(_2867_),
    .B1(_2945_),
    .B2(_2337_),
    .X(_2946_));
 sky130_fd_sc_hd__o211a_2 _6219_ (.A1(_2105_),
    .A2(_2802_),
    .B1(_2946_),
    .C1(_1085_),
    .X(_2947_));
 sky130_fd_sc_hd__o22a_2 _6220_ (.A1(_1060_),
    .A2(_2678_),
    .B1(_2737_),
    .B2(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__o22a_2 _6221_ (.A1(_2421_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(_2948_),
    .X(alu_out[28]));
 sky130_fd_sc_hd__o21ba_2 _6222_ (.A1(_1237_),
    .A2(_2741_),
    .B1_N(_2930_),
    .X(_2949_));
 sky130_fd_sc_hd__xnor2_2 _6223_ (.A(_1217_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__and2_2 _6224_ (.A(_1942_),
    .B(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__or2_2 _6225_ (.A(_1942_),
    .B(_2950_),
    .X(_2952_));
 sky130_fd_sc_hd__or2b_2 _6226_ (.A(_2951_),
    .B_N(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__a21oi_2 _6227_ (.A1(_2934_),
    .A2(_2940_),
    .B1(_2932_),
    .Y(_2954_));
 sky130_fd_sc_hd__or2_2 _6228_ (.A(_2953_),
    .B(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__nand2_2 _6229_ (.A(_2953_),
    .B(_2954_),
    .Y(_2956_));
 sky130_fd_sc_hd__and3_2 _6230_ (.A(_2503_),
    .B(_2955_),
    .C(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__or2b_2 _6231_ (.A(_2380_),
    .B_N(_2383_),
    .X(_2958_));
 sky130_fd_sc_hd__a21oi_2 _6232_ (.A1(_2923_),
    .A2(_2384_),
    .B1(_1148_),
    .Y(_2959_));
 sky130_fd_sc_hd__a211o_2 _6233_ (.A1(_1148_),
    .A2(_2958_),
    .B1(_2959_),
    .C1(_2337_),
    .X(_2960_));
 sky130_fd_sc_hd__o22a_2 _6234_ (.A1(_1111_),
    .A2(_2822_),
    .B1(_2896_),
    .B2(_2254_),
    .X(_2961_));
 sky130_fd_sc_hd__nor2_2 _6235_ (.A(_2102_),
    .B(_2692_),
    .Y(_2962_));
 sky130_fd_sc_hd__a32o_2 _6236_ (.A1(_1087_),
    .A2(_2960_),
    .A3(_2961_),
    .B1(_2962_),
    .B2(_1127_),
    .X(_2963_));
 sky130_fd_sc_hd__nor2_2 _6237_ (.A(_2701_),
    .B(_2797_),
    .Y(_2964_));
 sky130_fd_sc_hd__or3_2 _6238_ (.A(_2957_),
    .B(_2963_),
    .C(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__buf_1 _6239_ (.A(_2965_),
    .X(alu_out[29]));
 sky130_fd_sc_hd__or2_2 _6240_ (.A(_2442_),
    .B(_2942_),
    .X(_2966_));
 sky130_fd_sc_hd__inv_2 _6241_ (.A(_2547_),
    .Y(_2967_));
 sky130_fd_sc_hd__mux2_2 _6242_ (.A0(_2498_),
    .A1(_2967_),
    .S(_2327_),
    .X(_2968_));
 sky130_fd_sc_hd__mux2_2 _6243_ (.A0(_2420_),
    .A1(_2968_),
    .S(_2501_),
    .X(_2969_));
 sky130_fd_sc_hd__mux2_2 _6244_ (.A0(_2672_),
    .A1(_2674_),
    .S(_1803_),
    .X(_2970_));
 sky130_fd_sc_hd__mux2_2 _6245_ (.A0(_2675_),
    .A1(_2703_),
    .S(_1803_),
    .X(_2971_));
 sky130_fd_sc_hd__mux2_2 _6246_ (.A0(_2970_),
    .A1(_2971_),
    .S(_1126_),
    .X(_2972_));
 sky130_fd_sc_hd__inv_2 _6247_ (.A(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hd__mux2_2 _6248_ (.A0(_2969_),
    .A1(_2973_),
    .S(_2530_),
    .X(_2974_));
 sky130_fd_sc_hd__nand2_2 _6249_ (.A(_1148_),
    .B(_1925_),
    .Y(_2975_));
 sky130_fd_sc_hd__o31a_2 _6250_ (.A1(_2178_),
    .A2(_1980_),
    .A3(_1960_),
    .B1(_1127_),
    .X(_2976_));
 sky130_fd_sc_hd__o21ai_2 _6251_ (.A1(_1944_),
    .A2(_2975_),
    .B1(_2976_),
    .Y(_2977_));
 sky130_fd_sc_hd__o211a_2 _6252_ (.A1(_2104_),
    .A2(_2849_),
    .B1(_2977_),
    .C1(_1086_),
    .X(_2978_));
 sky130_fd_sc_hd__o21ai_2 _6253_ (.A1(_2255_),
    .A2(_2910_),
    .B1(_2978_),
    .Y(_2979_));
 sky130_fd_sc_hd__o211a_2 _6254_ (.A1(_2974_),
    .A2(_2797_),
    .B1(_2979_),
    .C1(_2421_),
    .X(_2980_));
 sky130_fd_sc_hd__nor2_2 _6255_ (.A(_1238_),
    .B(_2929_),
    .Y(_2981_));
 sky130_fd_sc_hd__nor2_2 _6256_ (.A(_2741_),
    .B(_2981_),
    .Y(_2982_));
 sky130_fd_sc_hd__xnor2_2 _6257_ (.A(_1348_),
    .B(_2982_),
    .Y(_2983_));
 sky130_fd_sc_hd__nor2_2 _6258_ (.A(_1923_),
    .B(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__and2_2 _6259_ (.A(_1923_),
    .B(_2983_),
    .X(_2985_));
 sky130_fd_sc_hd__nor2_2 _6260_ (.A(_2984_),
    .B(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__a211o_2 _6261_ (.A1(_2934_),
    .A2(_2940_),
    .B1(_2951_),
    .C1(_2932_),
    .X(_2987_));
 sky130_fd_sc_hd__and3_2 _6262_ (.A(_2952_),
    .B(_2986_),
    .C(_2987_),
    .X(_2988_));
 sky130_fd_sc_hd__a21oi_2 _6263_ (.A1(_2952_),
    .A2(_2987_),
    .B1(_2986_),
    .Y(_2989_));
 sky130_fd_sc_hd__nor2_2 _6264_ (.A(_2988_),
    .B(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__o2bb2a_2 _6265_ (.A1_N(_2966_),
    .A2_N(_2980_),
    .B1(_2408_),
    .B2(_2990_),
    .X(alu_out[30]));
 sky130_fd_sc_hd__a31o_2 _6266_ (.A1(_2952_),
    .A2(_2986_),
    .A3(_2987_),
    .B1(_2984_),
    .X(_2991_));
 sky130_fd_sc_hd__a21o_2 _6267_ (.A1(_1348_),
    .A2(_2981_),
    .B1(_2741_),
    .X(_2992_));
 sky130_fd_sc_hd__xor2_2 _6268_ (.A(_1334_),
    .B(_1904_),
    .X(_2993_));
 sky130_fd_sc_hd__xnor2_2 _6269_ (.A(_2992_),
    .B(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__xnor2_2 _6270_ (.A(_2991_),
    .B(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__inv_2 _6271_ (.A(_2942_),
    .Y(_2996_));
 sky130_fd_sc_hd__or2_2 _6272_ (.A(_2379_),
    .B(_2377_),
    .X(_2997_));
 sky130_fd_sc_hd__mux2_2 _6273_ (.A0(_2958_),
    .A1(_2997_),
    .S(_2363_),
    .X(_2998_));
 sky130_fd_sc_hd__o22a_2 _6274_ (.A1(_2254_),
    .A2(_2925_),
    .B1(_2998_),
    .B2(_2337_),
    .X(_2999_));
 sky130_fd_sc_hd__o211a_2 _6275_ (.A1(_2530_),
    .A2(_2859_),
    .B1(_2999_),
    .C1(_1087_),
    .X(_3000_));
 sky130_fd_sc_hd__a221o_2 _6276_ (.A1(_2720_),
    .A2(_2737_),
    .B1(_2996_),
    .B2(_2472_),
    .C1(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__o21bai_2 _6277_ (.A1(_2621_),
    .A2(_2995_),
    .B1_N(_3001_),
    .Y(alu_out[31]));
 sky130_fd_sc_hd__buf_1 _6278_ (.A(WD3[26]),
    .X(_3002_));
 sky130_fd_sc_hd__or3b_2 _6279_ (.A(A3[4]),
    .B(A3[2]),
    .C_N(A3[3]),
    .X(_3003_));
 sky130_fd_sc_hd__nand2_2 _6280_ (.A(A3[1]),
    .B(WE3),
    .Y(_3004_));
 sky130_fd_sc_hd__or2_2 _6281_ (.A(A3[0]),
    .B(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__nor2_2 _6282_ (.A(_3003_),
    .B(_3005_),
    .Y(_3006_));
 sky130_fd_sc_hd__buf_1 _6283_ (.A(_3006_),
    .X(_3007_));
 sky130_fd_sc_hd__mux2_2 _6284_ (.A0(\rf.registers[10][26] ),
    .A1(_3002_),
    .S(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__buf_1 _6285_ (.A(_3008_),
    .X(_0752_));
 sky130_fd_sc_hd__buf_1 _6286_ (.A(WD3[27]),
    .X(_3009_));
 sky130_fd_sc_hd__mux2_2 _6287_ (.A0(\rf.registers[10][27] ),
    .A1(_3009_),
    .S(_3007_),
    .X(_3010_));
 sky130_fd_sc_hd__buf_1 _6288_ (.A(_3010_),
    .X(_0753_));
 sky130_fd_sc_hd__buf_1 _6289_ (.A(WD3[28]),
    .X(_3011_));
 sky130_fd_sc_hd__mux2_2 _6290_ (.A0(\rf.registers[10][28] ),
    .A1(_3011_),
    .S(_3007_),
    .X(_3012_));
 sky130_fd_sc_hd__buf_1 _6291_ (.A(_3012_),
    .X(_0754_));
 sky130_fd_sc_hd__buf_1 _6292_ (.A(WD3[29]),
    .X(_3013_));
 sky130_fd_sc_hd__mux2_2 _6293_ (.A0(\rf.registers[10][29] ),
    .A1(_3013_),
    .S(_3007_),
    .X(_3014_));
 sky130_fd_sc_hd__buf_1 _6294_ (.A(_3014_),
    .X(_0755_));
 sky130_fd_sc_hd__buf_1 _6295_ (.A(WD3[30]),
    .X(_3015_));
 sky130_fd_sc_hd__mux2_2 _6296_ (.A0(\rf.registers[10][30] ),
    .A1(_3015_),
    .S(_3007_),
    .X(_3016_));
 sky130_fd_sc_hd__buf_1 _6297_ (.A(_3016_),
    .X(_0756_));
 sky130_fd_sc_hd__buf_1 _6298_ (.A(WD3[31]),
    .X(_3017_));
 sky130_fd_sc_hd__mux2_2 _6299_ (.A0(\rf.registers[10][31] ),
    .A1(_3017_),
    .S(_3007_),
    .X(_3018_));
 sky130_fd_sc_hd__buf_1 _6300_ (.A(_3018_),
    .X(_0757_));
 sky130_fd_sc_hd__buf_1 _6301_ (.A(WD3[0]),
    .X(_3019_));
 sky130_fd_sc_hd__nor2_2 _6302_ (.A(A3[0]),
    .B(_3004_),
    .Y(_3020_));
 sky130_fd_sc_hd__and3b_2 _6303_ (.A_N(A3[3]),
    .B(A3[2]),
    .C(A3[4]),
    .X(_3021_));
 sky130_fd_sc_hd__nand2_2 _6304_ (.A(_3020_),
    .B(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__buf_1 _6305_ (.A(_3022_),
    .X(_3023_));
 sky130_fd_sc_hd__mux2_2 _6306_ (.A0(_3019_),
    .A1(\rf.registers[22][0] ),
    .S(_3023_),
    .X(_3024_));
 sky130_fd_sc_hd__buf_1 _6307_ (.A(_3024_),
    .X(_0758_));
 sky130_fd_sc_hd__buf_1 _6308_ (.A(WD3[1]),
    .X(_3025_));
 sky130_fd_sc_hd__mux2_2 _6309_ (.A0(_3025_),
    .A1(\rf.registers[22][1] ),
    .S(_3023_),
    .X(_3026_));
 sky130_fd_sc_hd__buf_1 _6310_ (.A(_3026_),
    .X(_0759_));
 sky130_fd_sc_hd__buf_1 _6311_ (.A(WD3[2]),
    .X(_3027_));
 sky130_fd_sc_hd__mux2_2 _6312_ (.A0(_3027_),
    .A1(\rf.registers[22][2] ),
    .S(_3023_),
    .X(_3028_));
 sky130_fd_sc_hd__buf_1 _6313_ (.A(_3028_),
    .X(_0760_));
 sky130_fd_sc_hd__buf_1 _6314_ (.A(WD3[3]),
    .X(_3029_));
 sky130_fd_sc_hd__mux2_2 _6315_ (.A0(_3029_),
    .A1(\rf.registers[22][3] ),
    .S(_3023_),
    .X(_3030_));
 sky130_fd_sc_hd__buf_1 _6316_ (.A(_3030_),
    .X(_0761_));
 sky130_fd_sc_hd__buf_1 _6317_ (.A(WD3[4]),
    .X(_3031_));
 sky130_fd_sc_hd__mux2_2 _6318_ (.A0(_3031_),
    .A1(\rf.registers[22][4] ),
    .S(_3023_),
    .X(_3032_));
 sky130_fd_sc_hd__buf_1 _6319_ (.A(_3032_),
    .X(_0762_));
 sky130_fd_sc_hd__buf_1 _6320_ (.A(WD3[5]),
    .X(_3033_));
 sky130_fd_sc_hd__mux2_2 _6321_ (.A0(_3033_),
    .A1(\rf.registers[22][5] ),
    .S(_3023_),
    .X(_3034_));
 sky130_fd_sc_hd__buf_1 _6322_ (.A(_3034_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_1 _6323_ (.A(WD3[6]),
    .X(_3035_));
 sky130_fd_sc_hd__mux2_2 _6324_ (.A0(_3035_),
    .A1(\rf.registers[22][6] ),
    .S(_3023_),
    .X(_3036_));
 sky130_fd_sc_hd__buf_1 _6325_ (.A(_3036_),
    .X(_0764_));
 sky130_fd_sc_hd__buf_1 _6326_ (.A(WD3[7]),
    .X(_3037_));
 sky130_fd_sc_hd__mux2_2 _6327_ (.A0(_3037_),
    .A1(\rf.registers[22][7] ),
    .S(_3023_),
    .X(_3038_));
 sky130_fd_sc_hd__buf_1 _6328_ (.A(_3038_),
    .X(_0765_));
 sky130_fd_sc_hd__buf_1 _6329_ (.A(WD3[8]),
    .X(_3039_));
 sky130_fd_sc_hd__mux2_2 _6330_ (.A0(_3039_),
    .A1(\rf.registers[22][8] ),
    .S(_3023_),
    .X(_3040_));
 sky130_fd_sc_hd__buf_1 _6331_ (.A(_3040_),
    .X(_0766_));
 sky130_fd_sc_hd__buf_1 _6332_ (.A(WD3[9]),
    .X(_3041_));
 sky130_fd_sc_hd__mux2_2 _6333_ (.A0(_3041_),
    .A1(\rf.registers[22][9] ),
    .S(_3023_),
    .X(_3042_));
 sky130_fd_sc_hd__buf_1 _6334_ (.A(_3042_),
    .X(_0767_));
 sky130_fd_sc_hd__buf_1 _6335_ (.A(WD3[10]),
    .X(_3043_));
 sky130_fd_sc_hd__buf_1 _6336_ (.A(_3022_),
    .X(_3044_));
 sky130_fd_sc_hd__mux2_2 _6337_ (.A0(_3043_),
    .A1(\rf.registers[22][10] ),
    .S(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__buf_1 _6338_ (.A(_3045_),
    .X(_0768_));
 sky130_fd_sc_hd__buf_1 _6339_ (.A(WD3[11]),
    .X(_3046_));
 sky130_fd_sc_hd__mux2_2 _6340_ (.A0(_3046_),
    .A1(\rf.registers[22][11] ),
    .S(_3044_),
    .X(_3047_));
 sky130_fd_sc_hd__buf_1 _6341_ (.A(_3047_),
    .X(_0769_));
 sky130_fd_sc_hd__buf_1 _6342_ (.A(WD3[12]),
    .X(_3048_));
 sky130_fd_sc_hd__mux2_2 _6343_ (.A0(_3048_),
    .A1(\rf.registers[22][12] ),
    .S(_3044_),
    .X(_3049_));
 sky130_fd_sc_hd__buf_1 _6344_ (.A(_3049_),
    .X(_0770_));
 sky130_fd_sc_hd__buf_1 _6345_ (.A(WD3[13]),
    .X(_3050_));
 sky130_fd_sc_hd__mux2_2 _6346_ (.A0(_3050_),
    .A1(\rf.registers[22][13] ),
    .S(_3044_),
    .X(_3051_));
 sky130_fd_sc_hd__buf_1 _6347_ (.A(_3051_),
    .X(_0771_));
 sky130_fd_sc_hd__buf_1 _6348_ (.A(WD3[14]),
    .X(_3052_));
 sky130_fd_sc_hd__mux2_2 _6349_ (.A0(_3052_),
    .A1(\rf.registers[22][14] ),
    .S(_3044_),
    .X(_3053_));
 sky130_fd_sc_hd__buf_1 _6350_ (.A(_3053_),
    .X(_0772_));
 sky130_fd_sc_hd__buf_1 _6351_ (.A(WD3[15]),
    .X(_3054_));
 sky130_fd_sc_hd__mux2_2 _6352_ (.A0(_3054_),
    .A1(\rf.registers[22][15] ),
    .S(_3044_),
    .X(_3055_));
 sky130_fd_sc_hd__buf_1 _6353_ (.A(_3055_),
    .X(_0773_));
 sky130_fd_sc_hd__buf_1 _6354_ (.A(WD3[16]),
    .X(_3056_));
 sky130_fd_sc_hd__mux2_2 _6355_ (.A0(_3056_),
    .A1(\rf.registers[22][16] ),
    .S(_3044_),
    .X(_3057_));
 sky130_fd_sc_hd__buf_1 _6356_ (.A(_3057_),
    .X(_0774_));
 sky130_fd_sc_hd__buf_1 _6357_ (.A(WD3[17]),
    .X(_3058_));
 sky130_fd_sc_hd__mux2_2 _6358_ (.A0(_3058_),
    .A1(\rf.registers[22][17] ),
    .S(_3044_),
    .X(_3059_));
 sky130_fd_sc_hd__buf_1 _6359_ (.A(_3059_),
    .X(_0775_));
 sky130_fd_sc_hd__buf_1 _6360_ (.A(WD3[18]),
    .X(_3060_));
 sky130_fd_sc_hd__mux2_2 _6361_ (.A0(_3060_),
    .A1(\rf.registers[22][18] ),
    .S(_3044_),
    .X(_3061_));
 sky130_fd_sc_hd__buf_1 _6362_ (.A(_3061_),
    .X(_0776_));
 sky130_fd_sc_hd__buf_1 _6363_ (.A(WD3[19]),
    .X(_3062_));
 sky130_fd_sc_hd__mux2_2 _6364_ (.A0(_3062_),
    .A1(\rf.registers[22][19] ),
    .S(_3044_),
    .X(_3063_));
 sky130_fd_sc_hd__buf_1 _6365_ (.A(_3063_),
    .X(_0777_));
 sky130_fd_sc_hd__buf_1 _6366_ (.A(WD3[20]),
    .X(_3064_));
 sky130_fd_sc_hd__buf_1 _6367_ (.A(_3022_),
    .X(_3065_));
 sky130_fd_sc_hd__mux2_2 _6368_ (.A0(_3064_),
    .A1(\rf.registers[22][20] ),
    .S(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__buf_1 _6369_ (.A(_3066_),
    .X(_0778_));
 sky130_fd_sc_hd__buf_1 _6370_ (.A(WD3[21]),
    .X(_3067_));
 sky130_fd_sc_hd__mux2_2 _6371_ (.A0(_3067_),
    .A1(\rf.registers[22][21] ),
    .S(_3065_),
    .X(_3068_));
 sky130_fd_sc_hd__buf_1 _6372_ (.A(_3068_),
    .X(_0779_));
 sky130_fd_sc_hd__buf_1 _6373_ (.A(WD3[22]),
    .X(_3069_));
 sky130_fd_sc_hd__mux2_2 _6374_ (.A0(_3069_),
    .A1(\rf.registers[22][22] ),
    .S(_3065_),
    .X(_3070_));
 sky130_fd_sc_hd__buf_1 _6375_ (.A(_3070_),
    .X(_0780_));
 sky130_fd_sc_hd__buf_1 _6376_ (.A(WD3[23]),
    .X(_3071_));
 sky130_fd_sc_hd__mux2_2 _6377_ (.A0(_3071_),
    .A1(\rf.registers[22][23] ),
    .S(_3065_),
    .X(_3072_));
 sky130_fd_sc_hd__buf_1 _6378_ (.A(_3072_),
    .X(_0781_));
 sky130_fd_sc_hd__buf_1 _6379_ (.A(WD3[24]),
    .X(_3073_));
 sky130_fd_sc_hd__mux2_2 _6380_ (.A0(_3073_),
    .A1(\rf.registers[22][24] ),
    .S(_3065_),
    .X(_3074_));
 sky130_fd_sc_hd__buf_1 _6381_ (.A(_3074_),
    .X(_0782_));
 sky130_fd_sc_hd__buf_1 _6382_ (.A(WD3[25]),
    .X(_3075_));
 sky130_fd_sc_hd__mux2_2 _6383_ (.A0(_3075_),
    .A1(\rf.registers[22][25] ),
    .S(_3065_),
    .X(_3076_));
 sky130_fd_sc_hd__buf_1 _6384_ (.A(_3076_),
    .X(_0783_));
 sky130_fd_sc_hd__buf_1 _6385_ (.A(WD3[26]),
    .X(_3077_));
 sky130_fd_sc_hd__mux2_2 _6386_ (.A0(_3077_),
    .A1(\rf.registers[22][26] ),
    .S(_3065_),
    .X(_3078_));
 sky130_fd_sc_hd__buf_1 _6387_ (.A(_3078_),
    .X(_0784_));
 sky130_fd_sc_hd__buf_1 _6388_ (.A(WD3[27]),
    .X(_3079_));
 sky130_fd_sc_hd__mux2_2 _6389_ (.A0(_3079_),
    .A1(\rf.registers[22][27] ),
    .S(_3065_),
    .X(_3080_));
 sky130_fd_sc_hd__buf_1 _6390_ (.A(_3080_),
    .X(_0785_));
 sky130_fd_sc_hd__buf_1 _6391_ (.A(WD3[28]),
    .X(_3081_));
 sky130_fd_sc_hd__mux2_2 _6392_ (.A0(_3081_),
    .A1(\rf.registers[22][28] ),
    .S(_3065_),
    .X(_3082_));
 sky130_fd_sc_hd__buf_1 _6393_ (.A(_3082_),
    .X(_0786_));
 sky130_fd_sc_hd__buf_1 _6394_ (.A(WD3[29]),
    .X(_3083_));
 sky130_fd_sc_hd__mux2_2 _6395_ (.A0(_3083_),
    .A1(\rf.registers[22][29] ),
    .S(_3065_),
    .X(_3084_));
 sky130_fd_sc_hd__buf_1 _6396_ (.A(_3084_),
    .X(_0787_));
 sky130_fd_sc_hd__buf_1 _6397_ (.A(WD3[30]),
    .X(_3085_));
 sky130_fd_sc_hd__mux2_2 _6398_ (.A0(_3085_),
    .A1(\rf.registers[22][30] ),
    .S(_3022_),
    .X(_3086_));
 sky130_fd_sc_hd__buf_1 _6399_ (.A(_3086_),
    .X(_0788_));
 sky130_fd_sc_hd__buf_1 _6400_ (.A(WD3[31]),
    .X(_3087_));
 sky130_fd_sc_hd__mux2_2 _6401_ (.A0(_3087_),
    .A1(\rf.registers[22][31] ),
    .S(_3022_),
    .X(_3088_));
 sky130_fd_sc_hd__buf_1 _6402_ (.A(_3088_),
    .X(_0789_));
 sky130_fd_sc_hd__buf_1 _6403_ (.A(WD3[0]),
    .X(_3089_));
 sky130_fd_sc_hd__or3b_2 _6404_ (.A(A3[3]),
    .B(A3[2]),
    .C_N(A3[4]),
    .X(_3090_));
 sky130_fd_sc_hd__nand3b_2 _6405_ (.A_N(A3[1]),
    .B(A3[0]),
    .C(WE3),
    .Y(_3091_));
 sky130_fd_sc_hd__nor2_2 _6406_ (.A(_3090_),
    .B(_3091_),
    .Y(_3092_));
 sky130_fd_sc_hd__buf_1 _6407_ (.A(_3092_),
    .X(_3093_));
 sky130_fd_sc_hd__mux2_2 _6408_ (.A0(\rf.registers[17][0] ),
    .A1(_3089_),
    .S(_3093_),
    .X(_3094_));
 sky130_fd_sc_hd__buf_1 _6409_ (.A(_3094_),
    .X(_0790_));
 sky130_fd_sc_hd__buf_1 _6410_ (.A(WD3[1]),
    .X(_3095_));
 sky130_fd_sc_hd__mux2_2 _6411_ (.A0(\rf.registers[17][1] ),
    .A1(_3095_),
    .S(_3093_),
    .X(_3096_));
 sky130_fd_sc_hd__buf_1 _6412_ (.A(_3096_),
    .X(_0791_));
 sky130_fd_sc_hd__buf_1 _6413_ (.A(WD3[2]),
    .X(_3097_));
 sky130_fd_sc_hd__mux2_2 _6414_ (.A0(\rf.registers[17][2] ),
    .A1(_3097_),
    .S(_3093_),
    .X(_3098_));
 sky130_fd_sc_hd__buf_1 _6415_ (.A(_3098_),
    .X(_0792_));
 sky130_fd_sc_hd__buf_1 _6416_ (.A(WD3[3]),
    .X(_3099_));
 sky130_fd_sc_hd__mux2_2 _6417_ (.A0(\rf.registers[17][3] ),
    .A1(_3099_),
    .S(_3093_),
    .X(_3100_));
 sky130_fd_sc_hd__buf_1 _6418_ (.A(_3100_),
    .X(_0793_));
 sky130_fd_sc_hd__buf_1 _6419_ (.A(WD3[4]),
    .X(_3101_));
 sky130_fd_sc_hd__mux2_2 _6420_ (.A0(\rf.registers[17][4] ),
    .A1(_3101_),
    .S(_3093_),
    .X(_3102_));
 sky130_fd_sc_hd__buf_1 _6421_ (.A(_3102_),
    .X(_0794_));
 sky130_fd_sc_hd__buf_1 _6422_ (.A(WD3[5]),
    .X(_3103_));
 sky130_fd_sc_hd__mux2_2 _6423_ (.A0(\rf.registers[17][5] ),
    .A1(_3103_),
    .S(_3093_),
    .X(_3104_));
 sky130_fd_sc_hd__buf_1 _6424_ (.A(_3104_),
    .X(_0795_));
 sky130_fd_sc_hd__buf_1 _6425_ (.A(WD3[6]),
    .X(_3105_));
 sky130_fd_sc_hd__mux2_2 _6426_ (.A0(\rf.registers[17][6] ),
    .A1(_3105_),
    .S(_3093_),
    .X(_3106_));
 sky130_fd_sc_hd__buf_1 _6427_ (.A(_3106_),
    .X(_0796_));
 sky130_fd_sc_hd__buf_1 _6428_ (.A(WD3[7]),
    .X(_3107_));
 sky130_fd_sc_hd__mux2_2 _6429_ (.A0(\rf.registers[17][7] ),
    .A1(_3107_),
    .S(_3093_),
    .X(_3108_));
 sky130_fd_sc_hd__buf_1 _6430_ (.A(_3108_),
    .X(_0797_));
 sky130_fd_sc_hd__buf_1 _6431_ (.A(WD3[8]),
    .X(_3109_));
 sky130_fd_sc_hd__mux2_2 _6432_ (.A0(\rf.registers[17][8] ),
    .A1(_3109_),
    .S(_3093_),
    .X(_3110_));
 sky130_fd_sc_hd__buf_1 _6433_ (.A(_3110_),
    .X(_0798_));
 sky130_fd_sc_hd__buf_1 _6434_ (.A(WD3[9]),
    .X(_3111_));
 sky130_fd_sc_hd__mux2_2 _6435_ (.A0(\rf.registers[17][9] ),
    .A1(_3111_),
    .S(_3093_),
    .X(_3112_));
 sky130_fd_sc_hd__buf_1 _6436_ (.A(_3112_),
    .X(_0799_));
 sky130_fd_sc_hd__buf_1 _6437_ (.A(WD3[10]),
    .X(_3113_));
 sky130_fd_sc_hd__buf_1 _6438_ (.A(_3092_),
    .X(_3114_));
 sky130_fd_sc_hd__mux2_2 _6439_ (.A0(\rf.registers[17][10] ),
    .A1(_3113_),
    .S(_3114_),
    .X(_3115_));
 sky130_fd_sc_hd__buf_1 _6440_ (.A(_3115_),
    .X(_0800_));
 sky130_fd_sc_hd__buf_1 _6441_ (.A(WD3[11]),
    .X(_3116_));
 sky130_fd_sc_hd__mux2_2 _6442_ (.A0(\rf.registers[17][11] ),
    .A1(_3116_),
    .S(_3114_),
    .X(_3117_));
 sky130_fd_sc_hd__buf_1 _6443_ (.A(_3117_),
    .X(_0801_));
 sky130_fd_sc_hd__buf_1 _6444_ (.A(WD3[12]),
    .X(_3118_));
 sky130_fd_sc_hd__mux2_2 _6445_ (.A0(\rf.registers[17][12] ),
    .A1(_3118_),
    .S(_3114_),
    .X(_3119_));
 sky130_fd_sc_hd__buf_1 _6446_ (.A(_3119_),
    .X(_0802_));
 sky130_fd_sc_hd__buf_1 _6447_ (.A(WD3[13]),
    .X(_3120_));
 sky130_fd_sc_hd__mux2_2 _6448_ (.A0(\rf.registers[17][13] ),
    .A1(_3120_),
    .S(_3114_),
    .X(_3121_));
 sky130_fd_sc_hd__buf_1 _6449_ (.A(_3121_),
    .X(_0803_));
 sky130_fd_sc_hd__buf_1 _6450_ (.A(WD3[14]),
    .X(_3122_));
 sky130_fd_sc_hd__mux2_2 _6451_ (.A0(\rf.registers[17][14] ),
    .A1(_3122_),
    .S(_3114_),
    .X(_3123_));
 sky130_fd_sc_hd__buf_1 _6452_ (.A(_3123_),
    .X(_0804_));
 sky130_fd_sc_hd__buf_1 _6453_ (.A(WD3[15]),
    .X(_3124_));
 sky130_fd_sc_hd__mux2_2 _6454_ (.A0(\rf.registers[17][15] ),
    .A1(_3124_),
    .S(_3114_),
    .X(_3125_));
 sky130_fd_sc_hd__buf_1 _6455_ (.A(_3125_),
    .X(_0805_));
 sky130_fd_sc_hd__buf_1 _6456_ (.A(WD3[16]),
    .X(_3126_));
 sky130_fd_sc_hd__mux2_2 _6457_ (.A0(\rf.registers[17][16] ),
    .A1(_3126_),
    .S(_3114_),
    .X(_3127_));
 sky130_fd_sc_hd__buf_1 _6458_ (.A(_3127_),
    .X(_0806_));
 sky130_fd_sc_hd__buf_1 _6459_ (.A(WD3[17]),
    .X(_3128_));
 sky130_fd_sc_hd__mux2_2 _6460_ (.A0(\rf.registers[17][17] ),
    .A1(_3128_),
    .S(_3114_),
    .X(_3129_));
 sky130_fd_sc_hd__buf_1 _6461_ (.A(_3129_),
    .X(_0807_));
 sky130_fd_sc_hd__buf_1 _6462_ (.A(WD3[18]),
    .X(_3130_));
 sky130_fd_sc_hd__mux2_2 _6463_ (.A0(\rf.registers[17][18] ),
    .A1(_3130_),
    .S(_3114_),
    .X(_3131_));
 sky130_fd_sc_hd__buf_1 _6464_ (.A(_3131_),
    .X(_0808_));
 sky130_fd_sc_hd__buf_1 _6465_ (.A(WD3[19]),
    .X(_3132_));
 sky130_fd_sc_hd__mux2_2 _6466_ (.A0(\rf.registers[17][19] ),
    .A1(_3132_),
    .S(_3114_),
    .X(_3133_));
 sky130_fd_sc_hd__buf_1 _6467_ (.A(_3133_),
    .X(_0809_));
 sky130_fd_sc_hd__buf_1 _6468_ (.A(WD3[20]),
    .X(_3134_));
 sky130_fd_sc_hd__buf_1 _6469_ (.A(_3092_),
    .X(_3135_));
 sky130_fd_sc_hd__mux2_2 _6470_ (.A0(\rf.registers[17][20] ),
    .A1(_3134_),
    .S(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__buf_1 _6471_ (.A(_3136_),
    .X(_0810_));
 sky130_fd_sc_hd__buf_1 _6472_ (.A(WD3[21]),
    .X(_3137_));
 sky130_fd_sc_hd__mux2_2 _6473_ (.A0(\rf.registers[17][21] ),
    .A1(_3137_),
    .S(_3135_),
    .X(_3138_));
 sky130_fd_sc_hd__buf_1 _6474_ (.A(_3138_),
    .X(_0811_));
 sky130_fd_sc_hd__buf_1 _6475_ (.A(WD3[22]),
    .X(_3139_));
 sky130_fd_sc_hd__mux2_2 _6476_ (.A0(\rf.registers[17][22] ),
    .A1(_3139_),
    .S(_3135_),
    .X(_3140_));
 sky130_fd_sc_hd__buf_1 _6477_ (.A(_3140_),
    .X(_0812_));
 sky130_fd_sc_hd__buf_1 _6478_ (.A(WD3[23]),
    .X(_3141_));
 sky130_fd_sc_hd__mux2_2 _6479_ (.A0(\rf.registers[17][23] ),
    .A1(_3141_),
    .S(_3135_),
    .X(_3142_));
 sky130_fd_sc_hd__buf_1 _6480_ (.A(_3142_),
    .X(_0813_));
 sky130_fd_sc_hd__buf_1 _6481_ (.A(WD3[24]),
    .X(_3143_));
 sky130_fd_sc_hd__mux2_2 _6482_ (.A0(\rf.registers[17][24] ),
    .A1(_3143_),
    .S(_3135_),
    .X(_3144_));
 sky130_fd_sc_hd__buf_1 _6483_ (.A(_3144_),
    .X(_0814_));
 sky130_fd_sc_hd__buf_1 _6484_ (.A(WD3[25]),
    .X(_3145_));
 sky130_fd_sc_hd__mux2_2 _6485_ (.A0(\rf.registers[17][25] ),
    .A1(_3145_),
    .S(_3135_),
    .X(_3146_));
 sky130_fd_sc_hd__buf_1 _6486_ (.A(_3146_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_2 _6487_ (.A0(\rf.registers[17][26] ),
    .A1(_3002_),
    .S(_3135_),
    .X(_3147_));
 sky130_fd_sc_hd__buf_1 _6488_ (.A(_3147_),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_2 _6489_ (.A0(\rf.registers[17][27] ),
    .A1(_3009_),
    .S(_3135_),
    .X(_3148_));
 sky130_fd_sc_hd__buf_1 _6490_ (.A(_3148_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_2 _6491_ (.A0(\rf.registers[17][28] ),
    .A1(_3011_),
    .S(_3135_),
    .X(_3149_));
 sky130_fd_sc_hd__buf_1 _6492_ (.A(_3149_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_2 _6493_ (.A0(\rf.registers[17][29] ),
    .A1(_3013_),
    .S(_3135_),
    .X(_3150_));
 sky130_fd_sc_hd__buf_1 _6494_ (.A(_3150_),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_2 _6495_ (.A0(\rf.registers[17][30] ),
    .A1(_3015_),
    .S(_3092_),
    .X(_3151_));
 sky130_fd_sc_hd__buf_1 _6496_ (.A(_3151_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_2 _6497_ (.A0(\rf.registers[17][31] ),
    .A1(_3017_),
    .S(_3092_),
    .X(_3152_));
 sky130_fd_sc_hd__buf_1 _6498_ (.A(_3152_),
    .X(_0821_));
 sky130_fd_sc_hd__or3_2 _6499_ (.A(A3[4]),
    .B(A3[3]),
    .C(A3[2]),
    .X(_3153_));
 sky130_fd_sc_hd__or3b_2 _6500_ (.A(A3[1]),
    .B(A3[0]),
    .C_N(WE3),
    .X(_3154_));
 sky130_fd_sc_hd__buf_1 _6501_ (.A(_3154_),
    .X(_3155_));
 sky130_fd_sc_hd__nor2_2 _6502_ (.A(_3153_),
    .B(_3155_),
    .Y(_3156_));
 sky130_fd_sc_hd__buf_1 _6503_ (.A(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__mux2_2 _6504_ (.A0(\rf.registers[0][0] ),
    .A1(_3089_),
    .S(_3157_),
    .X(_3158_));
 sky130_fd_sc_hd__buf_1 _6505_ (.A(_3158_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_2 _6506_ (.A0(\rf.registers[0][1] ),
    .A1(_3095_),
    .S(_3157_),
    .X(_3159_));
 sky130_fd_sc_hd__buf_1 _6507_ (.A(_3159_),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_2 _6508_ (.A0(\rf.registers[0][2] ),
    .A1(_3097_),
    .S(_3157_),
    .X(_3160_));
 sky130_fd_sc_hd__buf_1 _6509_ (.A(_3160_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_2 _6510_ (.A0(\rf.registers[0][3] ),
    .A1(_3099_),
    .S(_3157_),
    .X(_3161_));
 sky130_fd_sc_hd__buf_1 _6511_ (.A(_3161_),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_2 _6512_ (.A0(\rf.registers[0][4] ),
    .A1(_3101_),
    .S(_3157_),
    .X(_3162_));
 sky130_fd_sc_hd__buf_1 _6513_ (.A(_3162_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_2 _6514_ (.A0(\rf.registers[0][5] ),
    .A1(_3103_),
    .S(_3157_),
    .X(_3163_));
 sky130_fd_sc_hd__buf_1 _6515_ (.A(_3163_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_2 _6516_ (.A0(\rf.registers[0][6] ),
    .A1(_3105_),
    .S(_3157_),
    .X(_3164_));
 sky130_fd_sc_hd__buf_1 _6517_ (.A(_3164_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_2 _6518_ (.A0(\rf.registers[0][7] ),
    .A1(_3107_),
    .S(_3157_),
    .X(_3165_));
 sky130_fd_sc_hd__buf_1 _6519_ (.A(_3165_),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_2 _6520_ (.A0(\rf.registers[0][8] ),
    .A1(_3109_),
    .S(_3157_),
    .X(_3166_));
 sky130_fd_sc_hd__buf_1 _6521_ (.A(_3166_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_2 _6522_ (.A0(\rf.registers[0][9] ),
    .A1(_3111_),
    .S(_3157_),
    .X(_3167_));
 sky130_fd_sc_hd__buf_1 _6523_ (.A(_3167_),
    .X(_0831_));
 sky130_fd_sc_hd__buf_1 _6524_ (.A(_3156_),
    .X(_3168_));
 sky130_fd_sc_hd__mux2_2 _6525_ (.A0(\rf.registers[0][10] ),
    .A1(_3113_),
    .S(_3168_),
    .X(_3169_));
 sky130_fd_sc_hd__buf_1 _6526_ (.A(_3169_),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_2 _6527_ (.A0(\rf.registers[0][11] ),
    .A1(_3116_),
    .S(_3168_),
    .X(_3170_));
 sky130_fd_sc_hd__buf_1 _6528_ (.A(_3170_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_2 _6529_ (.A0(\rf.registers[0][12] ),
    .A1(_3118_),
    .S(_3168_),
    .X(_3171_));
 sky130_fd_sc_hd__buf_1 _6530_ (.A(_3171_),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_2 _6531_ (.A0(\rf.registers[0][13] ),
    .A1(_3120_),
    .S(_3168_),
    .X(_3172_));
 sky130_fd_sc_hd__buf_1 _6532_ (.A(_3172_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_2 _6533_ (.A0(\rf.registers[0][14] ),
    .A1(_3122_),
    .S(_3168_),
    .X(_3173_));
 sky130_fd_sc_hd__buf_1 _6534_ (.A(_3173_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_2 _6535_ (.A0(\rf.registers[0][15] ),
    .A1(_3124_),
    .S(_3168_),
    .X(_3174_));
 sky130_fd_sc_hd__buf_1 _6536_ (.A(_3174_),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_2 _6537_ (.A0(\rf.registers[0][16] ),
    .A1(_3126_),
    .S(_3168_),
    .X(_3175_));
 sky130_fd_sc_hd__buf_1 _6538_ (.A(_3175_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_2 _6539_ (.A0(\rf.registers[0][17] ),
    .A1(_3128_),
    .S(_3168_),
    .X(_3176_));
 sky130_fd_sc_hd__buf_1 _6540_ (.A(_3176_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_2 _6541_ (.A0(\rf.registers[0][18] ),
    .A1(_3130_),
    .S(_3168_),
    .X(_3177_));
 sky130_fd_sc_hd__buf_1 _6542_ (.A(_3177_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_2 _6543_ (.A0(\rf.registers[0][19] ),
    .A1(_3132_),
    .S(_3168_),
    .X(_3178_));
 sky130_fd_sc_hd__buf_1 _6544_ (.A(_3178_),
    .X(_0841_));
 sky130_fd_sc_hd__buf_1 _6545_ (.A(_3156_),
    .X(_3179_));
 sky130_fd_sc_hd__mux2_2 _6546_ (.A0(\rf.registers[0][20] ),
    .A1(_3134_),
    .S(_3179_),
    .X(_3180_));
 sky130_fd_sc_hd__buf_1 _6547_ (.A(_3180_),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_2 _6548_ (.A0(\rf.registers[0][21] ),
    .A1(_3137_),
    .S(_3179_),
    .X(_3181_));
 sky130_fd_sc_hd__buf_1 _6549_ (.A(_3181_),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_2 _6550_ (.A0(\rf.registers[0][22] ),
    .A1(_3139_),
    .S(_3179_),
    .X(_3182_));
 sky130_fd_sc_hd__buf_1 _6551_ (.A(_3182_),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_2 _6552_ (.A0(\rf.registers[0][23] ),
    .A1(_3141_),
    .S(_3179_),
    .X(_3183_));
 sky130_fd_sc_hd__buf_1 _6553_ (.A(_3183_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_2 _6554_ (.A0(\rf.registers[0][24] ),
    .A1(_3143_),
    .S(_3179_),
    .X(_3184_));
 sky130_fd_sc_hd__buf_1 _6555_ (.A(_3184_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_2 _6556_ (.A0(\rf.registers[0][25] ),
    .A1(_3145_),
    .S(_3179_),
    .X(_3185_));
 sky130_fd_sc_hd__buf_1 _6557_ (.A(_3185_),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_2 _6558_ (.A0(\rf.registers[0][26] ),
    .A1(_3002_),
    .S(_3179_),
    .X(_3186_));
 sky130_fd_sc_hd__buf_1 _6559_ (.A(_3186_),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_2 _6560_ (.A0(\rf.registers[0][27] ),
    .A1(_3009_),
    .S(_3179_),
    .X(_3187_));
 sky130_fd_sc_hd__buf_1 _6561_ (.A(_3187_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_2 _6562_ (.A0(\rf.registers[0][28] ),
    .A1(_3011_),
    .S(_3179_),
    .X(_3188_));
 sky130_fd_sc_hd__buf_1 _6563_ (.A(_3188_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_2 _6564_ (.A0(\rf.registers[0][29] ),
    .A1(_3013_),
    .S(_3179_),
    .X(_3189_));
 sky130_fd_sc_hd__buf_1 _6565_ (.A(_3189_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_2 _6566_ (.A0(\rf.registers[0][30] ),
    .A1(_3015_),
    .S(_3156_),
    .X(_3190_));
 sky130_fd_sc_hd__buf_1 _6567_ (.A(_3190_),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_2 _6568_ (.A0(\rf.registers[0][31] ),
    .A1(_3017_),
    .S(_3156_),
    .X(_3191_));
 sky130_fd_sc_hd__buf_1 _6569_ (.A(_3191_),
    .X(_0853_));
 sky130_fd_sc_hd__and3b_2 _6570_ (.A_N(A3[4]),
    .B(A3[3]),
    .C(A3[2]),
    .X(_3192_));
 sky130_fd_sc_hd__and3_2 _6571_ (.A(A3[1]),
    .B(A3[0]),
    .C(WE3),
    .X(_3193_));
 sky130_fd_sc_hd__nand2_2 _6572_ (.A(_3192_),
    .B(_3193_),
    .Y(_3194_));
 sky130_fd_sc_hd__buf_1 _6573_ (.A(_3194_),
    .X(_3195_));
 sky130_fd_sc_hd__mux2_2 _6574_ (.A0(_3019_),
    .A1(\rf.registers[15][0] ),
    .S(_3195_),
    .X(_3196_));
 sky130_fd_sc_hd__buf_1 _6575_ (.A(_3196_),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_2 _6576_ (.A0(_3025_),
    .A1(\rf.registers[15][1] ),
    .S(_3195_),
    .X(_3197_));
 sky130_fd_sc_hd__buf_1 _6577_ (.A(_3197_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_2 _6578_ (.A0(_3027_),
    .A1(\rf.registers[15][2] ),
    .S(_3195_),
    .X(_3198_));
 sky130_fd_sc_hd__buf_1 _6579_ (.A(_3198_),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_2 _6580_ (.A0(_3029_),
    .A1(\rf.registers[15][3] ),
    .S(_3195_),
    .X(_3199_));
 sky130_fd_sc_hd__buf_1 _6581_ (.A(_3199_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_2 _6582_ (.A0(_3031_),
    .A1(\rf.registers[15][4] ),
    .S(_3195_),
    .X(_3200_));
 sky130_fd_sc_hd__buf_1 _6583_ (.A(_3200_),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_2 _6584_ (.A0(_3033_),
    .A1(\rf.registers[15][5] ),
    .S(_3195_),
    .X(_3201_));
 sky130_fd_sc_hd__buf_1 _6585_ (.A(_3201_),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_2 _6586_ (.A0(_3035_),
    .A1(\rf.registers[15][6] ),
    .S(_3195_),
    .X(_3202_));
 sky130_fd_sc_hd__buf_1 _6587_ (.A(_3202_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_2 _6588_ (.A0(_3037_),
    .A1(\rf.registers[15][7] ),
    .S(_3195_),
    .X(_3203_));
 sky130_fd_sc_hd__buf_1 _6589_ (.A(_3203_),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_2 _6590_ (.A0(_3039_),
    .A1(\rf.registers[15][8] ),
    .S(_3195_),
    .X(_3204_));
 sky130_fd_sc_hd__buf_1 _6591_ (.A(_3204_),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_2 _6592_ (.A0(_3041_),
    .A1(\rf.registers[15][9] ),
    .S(_3195_),
    .X(_3205_));
 sky130_fd_sc_hd__buf_1 _6593_ (.A(_3205_),
    .X(_0863_));
 sky130_fd_sc_hd__buf_1 _6594_ (.A(_3194_),
    .X(_3206_));
 sky130_fd_sc_hd__mux2_2 _6595_ (.A0(_3043_),
    .A1(\rf.registers[15][10] ),
    .S(_3206_),
    .X(_3207_));
 sky130_fd_sc_hd__buf_1 _6596_ (.A(_3207_),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_2 _6597_ (.A0(_3046_),
    .A1(\rf.registers[15][11] ),
    .S(_3206_),
    .X(_3208_));
 sky130_fd_sc_hd__buf_1 _6598_ (.A(_3208_),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_2 _6599_ (.A0(_3048_),
    .A1(\rf.registers[15][12] ),
    .S(_3206_),
    .X(_3209_));
 sky130_fd_sc_hd__buf_1 _6600_ (.A(_3209_),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_2 _6601_ (.A0(_3050_),
    .A1(\rf.registers[15][13] ),
    .S(_3206_),
    .X(_3210_));
 sky130_fd_sc_hd__buf_1 _6602_ (.A(_3210_),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_2 _6603_ (.A0(_3052_),
    .A1(\rf.registers[15][14] ),
    .S(_3206_),
    .X(_3211_));
 sky130_fd_sc_hd__buf_1 _6604_ (.A(_3211_),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_2 _6605_ (.A0(_3054_),
    .A1(\rf.registers[15][15] ),
    .S(_3206_),
    .X(_3212_));
 sky130_fd_sc_hd__buf_1 _6606_ (.A(_3212_),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_2 _6607_ (.A0(_3056_),
    .A1(\rf.registers[15][16] ),
    .S(_3206_),
    .X(_3213_));
 sky130_fd_sc_hd__buf_1 _6608_ (.A(_3213_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_2 _6609_ (.A0(_3058_),
    .A1(\rf.registers[15][17] ),
    .S(_3206_),
    .X(_3214_));
 sky130_fd_sc_hd__buf_1 _6610_ (.A(_3214_),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_2 _6611_ (.A0(_3060_),
    .A1(\rf.registers[15][18] ),
    .S(_3206_),
    .X(_3215_));
 sky130_fd_sc_hd__buf_1 _6612_ (.A(_3215_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_2 _6613_ (.A0(_3062_),
    .A1(\rf.registers[15][19] ),
    .S(_3206_),
    .X(_3216_));
 sky130_fd_sc_hd__buf_1 _6614_ (.A(_3216_),
    .X(_0873_));
 sky130_fd_sc_hd__buf_1 _6615_ (.A(_3194_),
    .X(_3217_));
 sky130_fd_sc_hd__mux2_2 _6616_ (.A0(_3064_),
    .A1(\rf.registers[15][20] ),
    .S(_3217_),
    .X(_3218_));
 sky130_fd_sc_hd__buf_1 _6617_ (.A(_3218_),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_2 _6618_ (.A0(_3067_),
    .A1(\rf.registers[15][21] ),
    .S(_3217_),
    .X(_3219_));
 sky130_fd_sc_hd__buf_1 _6619_ (.A(_3219_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_2 _6620_ (.A0(_3069_),
    .A1(\rf.registers[15][22] ),
    .S(_3217_),
    .X(_3220_));
 sky130_fd_sc_hd__buf_1 _6621_ (.A(_3220_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_2 _6622_ (.A0(_3071_),
    .A1(\rf.registers[15][23] ),
    .S(_3217_),
    .X(_3221_));
 sky130_fd_sc_hd__buf_1 _6623_ (.A(_3221_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_2 _6624_ (.A0(_3073_),
    .A1(\rf.registers[15][24] ),
    .S(_3217_),
    .X(_3222_));
 sky130_fd_sc_hd__buf_1 _6625_ (.A(_3222_),
    .X(_0878_));
 sky130_fd_sc_hd__mux2_2 _6626_ (.A0(_3075_),
    .A1(\rf.registers[15][25] ),
    .S(_3217_),
    .X(_3223_));
 sky130_fd_sc_hd__buf_1 _6627_ (.A(_3223_),
    .X(_0879_));
 sky130_fd_sc_hd__mux2_2 _6628_ (.A0(_3077_),
    .A1(\rf.registers[15][26] ),
    .S(_3217_),
    .X(_3224_));
 sky130_fd_sc_hd__buf_1 _6629_ (.A(_3224_),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_2 _6630_ (.A0(_3079_),
    .A1(\rf.registers[15][27] ),
    .S(_3217_),
    .X(_3225_));
 sky130_fd_sc_hd__buf_1 _6631_ (.A(_3225_),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_2 _6632_ (.A0(_3081_),
    .A1(\rf.registers[15][28] ),
    .S(_3217_),
    .X(_3226_));
 sky130_fd_sc_hd__buf_1 _6633_ (.A(_3226_),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_2 _6634_ (.A0(_3083_),
    .A1(\rf.registers[15][29] ),
    .S(_3217_),
    .X(_3227_));
 sky130_fd_sc_hd__buf_1 _6635_ (.A(_3227_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_2 _6636_ (.A0(_3085_),
    .A1(\rf.registers[15][30] ),
    .S(_3194_),
    .X(_3228_));
 sky130_fd_sc_hd__buf_1 _6637_ (.A(_3228_),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_2 _6638_ (.A0(_3087_),
    .A1(\rf.registers[15][31] ),
    .S(_3194_),
    .X(_3229_));
 sky130_fd_sc_hd__buf_1 _6639_ (.A(_3229_),
    .X(_0885_));
 sky130_fd_sc_hd__nor2_2 _6640_ (.A(_3003_),
    .B(_3155_),
    .Y(_3230_));
 sky130_fd_sc_hd__buf_1 _6641_ (.A(_3230_),
    .X(_3231_));
 sky130_fd_sc_hd__mux2_2 _6642_ (.A0(\rf.registers[8][0] ),
    .A1(_3089_),
    .S(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__buf_1 _6643_ (.A(_3232_),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_2 _6644_ (.A0(\rf.registers[8][1] ),
    .A1(_3095_),
    .S(_3231_),
    .X(_3233_));
 sky130_fd_sc_hd__buf_1 _6645_ (.A(_3233_),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_2 _6646_ (.A0(\rf.registers[8][2] ),
    .A1(_3097_),
    .S(_3231_),
    .X(_3234_));
 sky130_fd_sc_hd__buf_1 _6647_ (.A(_3234_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_2 _6648_ (.A0(\rf.registers[8][3] ),
    .A1(_3099_),
    .S(_3231_),
    .X(_3235_));
 sky130_fd_sc_hd__buf_1 _6649_ (.A(_3235_),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_2 _6650_ (.A0(\rf.registers[8][4] ),
    .A1(_3101_),
    .S(_3231_),
    .X(_3236_));
 sky130_fd_sc_hd__buf_1 _6651_ (.A(_3236_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_2 _6652_ (.A0(\rf.registers[8][5] ),
    .A1(_3103_),
    .S(_3231_),
    .X(_3237_));
 sky130_fd_sc_hd__buf_1 _6653_ (.A(_3237_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_2 _6654_ (.A0(\rf.registers[8][6] ),
    .A1(_3105_),
    .S(_3231_),
    .X(_3238_));
 sky130_fd_sc_hd__buf_1 _6655_ (.A(_3238_),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_2 _6656_ (.A0(\rf.registers[8][7] ),
    .A1(_3107_),
    .S(_3231_),
    .X(_3239_));
 sky130_fd_sc_hd__buf_1 _6657_ (.A(_3239_),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_2 _6658_ (.A0(\rf.registers[8][8] ),
    .A1(_3109_),
    .S(_3231_),
    .X(_3240_));
 sky130_fd_sc_hd__buf_1 _6659_ (.A(_3240_),
    .X(_0894_));
 sky130_fd_sc_hd__mux2_2 _6660_ (.A0(\rf.registers[8][9] ),
    .A1(_3111_),
    .S(_3231_),
    .X(_3241_));
 sky130_fd_sc_hd__buf_1 _6661_ (.A(_3241_),
    .X(_0895_));
 sky130_fd_sc_hd__buf_1 _6662_ (.A(_3230_),
    .X(_3242_));
 sky130_fd_sc_hd__mux2_2 _6663_ (.A0(\rf.registers[8][10] ),
    .A1(_3113_),
    .S(_3242_),
    .X(_3243_));
 sky130_fd_sc_hd__buf_1 _6664_ (.A(_3243_),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_2 _6665_ (.A0(\rf.registers[8][11] ),
    .A1(_3116_),
    .S(_3242_),
    .X(_3244_));
 sky130_fd_sc_hd__buf_1 _6666_ (.A(_3244_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_2 _6667_ (.A0(\rf.registers[8][12] ),
    .A1(_3118_),
    .S(_3242_),
    .X(_3245_));
 sky130_fd_sc_hd__buf_1 _6668_ (.A(_3245_),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_2 _6669_ (.A0(\rf.registers[8][13] ),
    .A1(_3120_),
    .S(_3242_),
    .X(_3246_));
 sky130_fd_sc_hd__buf_1 _6670_ (.A(_3246_),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_2 _6671_ (.A0(\rf.registers[8][14] ),
    .A1(_3122_),
    .S(_3242_),
    .X(_3247_));
 sky130_fd_sc_hd__buf_1 _6672_ (.A(_3247_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_2 _6673_ (.A0(\rf.registers[8][15] ),
    .A1(_3124_),
    .S(_3242_),
    .X(_3248_));
 sky130_fd_sc_hd__buf_1 _6674_ (.A(_3248_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_2 _6675_ (.A0(\rf.registers[8][16] ),
    .A1(_3126_),
    .S(_3242_),
    .X(_3249_));
 sky130_fd_sc_hd__buf_1 _6676_ (.A(_3249_),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_2 _6677_ (.A0(\rf.registers[8][17] ),
    .A1(_3128_),
    .S(_3242_),
    .X(_3250_));
 sky130_fd_sc_hd__buf_1 _6678_ (.A(_3250_),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_2 _6679_ (.A0(\rf.registers[8][18] ),
    .A1(_3130_),
    .S(_3242_),
    .X(_3251_));
 sky130_fd_sc_hd__buf_1 _6680_ (.A(_3251_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_2 _6681_ (.A0(\rf.registers[8][19] ),
    .A1(_3132_),
    .S(_3242_),
    .X(_3252_));
 sky130_fd_sc_hd__buf_1 _6682_ (.A(_3252_),
    .X(_0905_));
 sky130_fd_sc_hd__buf_1 _6683_ (.A(_3230_),
    .X(_3253_));
 sky130_fd_sc_hd__mux2_2 _6684_ (.A0(\rf.registers[8][20] ),
    .A1(_3134_),
    .S(_3253_),
    .X(_3254_));
 sky130_fd_sc_hd__buf_1 _6685_ (.A(_3254_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_2 _6686_ (.A0(\rf.registers[8][21] ),
    .A1(_3137_),
    .S(_3253_),
    .X(_3255_));
 sky130_fd_sc_hd__buf_1 _6687_ (.A(_3255_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_2 _6688_ (.A0(\rf.registers[8][22] ),
    .A1(_3139_),
    .S(_3253_),
    .X(_3256_));
 sky130_fd_sc_hd__buf_1 _6689_ (.A(_3256_),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_2 _6690_ (.A0(\rf.registers[8][23] ),
    .A1(_3141_),
    .S(_3253_),
    .X(_3257_));
 sky130_fd_sc_hd__buf_1 _6691_ (.A(_3257_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_2 _6692_ (.A0(\rf.registers[8][24] ),
    .A1(_3143_),
    .S(_3253_),
    .X(_3258_));
 sky130_fd_sc_hd__buf_1 _6693_ (.A(_3258_),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_2 _6694_ (.A0(\rf.registers[8][25] ),
    .A1(_3145_),
    .S(_3253_),
    .X(_3259_));
 sky130_fd_sc_hd__buf_1 _6695_ (.A(_3259_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_2 _6696_ (.A0(\rf.registers[8][26] ),
    .A1(_3002_),
    .S(_3253_),
    .X(_3260_));
 sky130_fd_sc_hd__buf_1 _6697_ (.A(_3260_),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_2 _6698_ (.A0(\rf.registers[8][27] ),
    .A1(_3009_),
    .S(_3253_),
    .X(_3261_));
 sky130_fd_sc_hd__buf_1 _6699_ (.A(_3261_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_2 _6700_ (.A0(\rf.registers[8][28] ),
    .A1(_3011_),
    .S(_3253_),
    .X(_3262_));
 sky130_fd_sc_hd__buf_1 _6701_ (.A(_3262_),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_2 _6702_ (.A0(\rf.registers[8][29] ),
    .A1(_3013_),
    .S(_3253_),
    .X(_3263_));
 sky130_fd_sc_hd__buf_1 _6703_ (.A(_3263_),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_2 _6704_ (.A0(\rf.registers[8][30] ),
    .A1(_3015_),
    .S(_3230_),
    .X(_3264_));
 sky130_fd_sc_hd__buf_1 _6705_ (.A(_3264_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_2 _6706_ (.A0(\rf.registers[8][31] ),
    .A1(_3017_),
    .S(_3230_),
    .X(_3265_));
 sky130_fd_sc_hd__buf_1 _6707_ (.A(_3265_),
    .X(_0917_));
 sky130_fd_sc_hd__nand2_2 _6708_ (.A(_3020_),
    .B(_3192_),
    .Y(_3266_));
 sky130_fd_sc_hd__buf_1 _6709_ (.A(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__mux2_2 _6710_ (.A0(_3019_),
    .A1(\rf.registers[14][0] ),
    .S(_3267_),
    .X(_3268_));
 sky130_fd_sc_hd__buf_1 _6711_ (.A(_3268_),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_2 _6712_ (.A0(_3025_),
    .A1(\rf.registers[14][1] ),
    .S(_3267_),
    .X(_3269_));
 sky130_fd_sc_hd__buf_1 _6713_ (.A(_3269_),
    .X(_0919_));
 sky130_fd_sc_hd__mux2_2 _6714_ (.A0(_3027_),
    .A1(\rf.registers[14][2] ),
    .S(_3267_),
    .X(_3270_));
 sky130_fd_sc_hd__buf_1 _6715_ (.A(_3270_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_2 _6716_ (.A0(_3029_),
    .A1(\rf.registers[14][3] ),
    .S(_3267_),
    .X(_3271_));
 sky130_fd_sc_hd__buf_1 _6717_ (.A(_3271_),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_2 _6718_ (.A0(_3031_),
    .A1(\rf.registers[14][4] ),
    .S(_3267_),
    .X(_3272_));
 sky130_fd_sc_hd__buf_1 _6719_ (.A(_3272_),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_2 _6720_ (.A0(_3033_),
    .A1(\rf.registers[14][5] ),
    .S(_3267_),
    .X(_3273_));
 sky130_fd_sc_hd__buf_1 _6721_ (.A(_3273_),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_2 _6722_ (.A0(_3035_),
    .A1(\rf.registers[14][6] ),
    .S(_3267_),
    .X(_3274_));
 sky130_fd_sc_hd__buf_1 _6723_ (.A(_3274_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_2 _6724_ (.A0(_3037_),
    .A1(\rf.registers[14][7] ),
    .S(_3267_),
    .X(_3275_));
 sky130_fd_sc_hd__buf_1 _6725_ (.A(_3275_),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_2 _6726_ (.A0(_3039_),
    .A1(\rf.registers[14][8] ),
    .S(_3267_),
    .X(_3276_));
 sky130_fd_sc_hd__buf_1 _6727_ (.A(_3276_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_2 _6728_ (.A0(_3041_),
    .A1(\rf.registers[14][9] ),
    .S(_3267_),
    .X(_3277_));
 sky130_fd_sc_hd__buf_1 _6729_ (.A(_3277_),
    .X(_0927_));
 sky130_fd_sc_hd__buf_1 _6730_ (.A(_3266_),
    .X(_3278_));
 sky130_fd_sc_hd__mux2_2 _6731_ (.A0(_3043_),
    .A1(\rf.registers[14][10] ),
    .S(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__buf_1 _6732_ (.A(_3279_),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_2 _6733_ (.A0(_3046_),
    .A1(\rf.registers[14][11] ),
    .S(_3278_),
    .X(_3280_));
 sky130_fd_sc_hd__buf_1 _6734_ (.A(_3280_),
    .X(_0929_));
 sky130_fd_sc_hd__mux2_2 _6735_ (.A0(_3048_),
    .A1(\rf.registers[14][12] ),
    .S(_3278_),
    .X(_3281_));
 sky130_fd_sc_hd__buf_1 _6736_ (.A(_3281_),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_2 _6737_ (.A0(_3050_),
    .A1(\rf.registers[14][13] ),
    .S(_3278_),
    .X(_3282_));
 sky130_fd_sc_hd__buf_1 _6738_ (.A(_3282_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_2 _6739_ (.A0(_3052_),
    .A1(\rf.registers[14][14] ),
    .S(_3278_),
    .X(_3283_));
 sky130_fd_sc_hd__buf_1 _6740_ (.A(_3283_),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_2 _6741_ (.A0(_3054_),
    .A1(\rf.registers[14][15] ),
    .S(_3278_),
    .X(_3284_));
 sky130_fd_sc_hd__buf_1 _6742_ (.A(_3284_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_2 _6743_ (.A0(_3056_),
    .A1(\rf.registers[14][16] ),
    .S(_3278_),
    .X(_3285_));
 sky130_fd_sc_hd__buf_1 _6744_ (.A(_3285_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_2 _6745_ (.A0(_3058_),
    .A1(\rf.registers[14][17] ),
    .S(_3278_),
    .X(_3286_));
 sky130_fd_sc_hd__buf_1 _6746_ (.A(_3286_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_2 _6747_ (.A0(_3060_),
    .A1(\rf.registers[14][18] ),
    .S(_3278_),
    .X(_3287_));
 sky130_fd_sc_hd__buf_1 _6748_ (.A(_3287_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_2 _6749_ (.A0(_3062_),
    .A1(\rf.registers[14][19] ),
    .S(_3278_),
    .X(_3288_));
 sky130_fd_sc_hd__buf_1 _6750_ (.A(_3288_),
    .X(_0937_));
 sky130_fd_sc_hd__buf_1 _6751_ (.A(_3266_),
    .X(_3289_));
 sky130_fd_sc_hd__mux2_2 _6752_ (.A0(_3064_),
    .A1(\rf.registers[14][20] ),
    .S(_3289_),
    .X(_3290_));
 sky130_fd_sc_hd__buf_1 _6753_ (.A(_3290_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_2 _6754_ (.A0(_3067_),
    .A1(\rf.registers[14][21] ),
    .S(_3289_),
    .X(_3291_));
 sky130_fd_sc_hd__buf_1 _6755_ (.A(_3291_),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_2 _6756_ (.A0(_3069_),
    .A1(\rf.registers[14][22] ),
    .S(_3289_),
    .X(_3292_));
 sky130_fd_sc_hd__buf_1 _6757_ (.A(_3292_),
    .X(_0940_));
 sky130_fd_sc_hd__mux2_2 _6758_ (.A0(_3071_),
    .A1(\rf.registers[14][23] ),
    .S(_3289_),
    .X(_3293_));
 sky130_fd_sc_hd__buf_1 _6759_ (.A(_3293_),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_2 _6760_ (.A0(_3073_),
    .A1(\rf.registers[14][24] ),
    .S(_3289_),
    .X(_3294_));
 sky130_fd_sc_hd__buf_1 _6761_ (.A(_3294_),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_2 _6762_ (.A0(_3075_),
    .A1(\rf.registers[14][25] ),
    .S(_3289_),
    .X(_3295_));
 sky130_fd_sc_hd__buf_1 _6763_ (.A(_3295_),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_2 _6764_ (.A0(_3077_),
    .A1(\rf.registers[14][26] ),
    .S(_3289_),
    .X(_3296_));
 sky130_fd_sc_hd__buf_1 _6765_ (.A(_3296_),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_2 _6766_ (.A0(_3079_),
    .A1(\rf.registers[14][27] ),
    .S(_3289_),
    .X(_3297_));
 sky130_fd_sc_hd__buf_1 _6767_ (.A(_3297_),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_2 _6768_ (.A0(_3081_),
    .A1(\rf.registers[14][28] ),
    .S(_3289_),
    .X(_3298_));
 sky130_fd_sc_hd__buf_1 _6769_ (.A(_3298_),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_2 _6770_ (.A0(_3083_),
    .A1(\rf.registers[14][29] ),
    .S(_3289_),
    .X(_3299_));
 sky130_fd_sc_hd__buf_1 _6771_ (.A(_3299_),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_2 _6772_ (.A0(_3085_),
    .A1(\rf.registers[14][30] ),
    .S(_3266_),
    .X(_3300_));
 sky130_fd_sc_hd__buf_1 _6773_ (.A(_3300_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_2 _6774_ (.A0(_3087_),
    .A1(\rf.registers[14][31] ),
    .S(_3266_),
    .X(_3301_));
 sky130_fd_sc_hd__buf_1 _6775_ (.A(_3301_),
    .X(_0949_));
 sky130_fd_sc_hd__or3b_2 _6776_ (.A(A3[4]),
    .B(A3[3]),
    .C_N(A3[2]),
    .X(_3302_));
 sky130_fd_sc_hd__nor2_2 _6777_ (.A(_3005_),
    .B(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__buf_1 _6778_ (.A(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__mux2_2 _6779_ (.A0(\rf.registers[6][0] ),
    .A1(_3089_),
    .S(_3304_),
    .X(_3305_));
 sky130_fd_sc_hd__buf_1 _6780_ (.A(_3305_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_2 _6781_ (.A0(\rf.registers[6][1] ),
    .A1(_3095_),
    .S(_3304_),
    .X(_3306_));
 sky130_fd_sc_hd__buf_1 _6782_ (.A(_3306_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_2 _6783_ (.A0(\rf.registers[6][2] ),
    .A1(_3097_),
    .S(_3304_),
    .X(_3307_));
 sky130_fd_sc_hd__buf_1 _6784_ (.A(_3307_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_2 _6785_ (.A0(\rf.registers[6][3] ),
    .A1(_3099_),
    .S(_3304_),
    .X(_3308_));
 sky130_fd_sc_hd__buf_1 _6786_ (.A(_3308_),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_2 _6787_ (.A0(\rf.registers[6][4] ),
    .A1(_3101_),
    .S(_3304_),
    .X(_3309_));
 sky130_fd_sc_hd__buf_1 _6788_ (.A(_3309_),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_2 _6789_ (.A0(\rf.registers[6][5] ),
    .A1(_3103_),
    .S(_3304_),
    .X(_3310_));
 sky130_fd_sc_hd__buf_1 _6790_ (.A(_3310_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_2 _6791_ (.A0(\rf.registers[6][6] ),
    .A1(_3105_),
    .S(_3304_),
    .X(_3311_));
 sky130_fd_sc_hd__buf_1 _6792_ (.A(_3311_),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_2 _6793_ (.A0(\rf.registers[6][7] ),
    .A1(_3107_),
    .S(_3304_),
    .X(_3312_));
 sky130_fd_sc_hd__buf_1 _6794_ (.A(_3312_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_2 _6795_ (.A0(\rf.registers[6][8] ),
    .A1(_3109_),
    .S(_3304_),
    .X(_3313_));
 sky130_fd_sc_hd__buf_1 _6796_ (.A(_3313_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_2 _6797_ (.A0(\rf.registers[6][9] ),
    .A1(_3111_),
    .S(_3304_),
    .X(_3314_));
 sky130_fd_sc_hd__buf_1 _6798_ (.A(_3314_),
    .X(_0959_));
 sky130_fd_sc_hd__buf_1 _6799_ (.A(_3303_),
    .X(_3315_));
 sky130_fd_sc_hd__mux2_2 _6800_ (.A0(\rf.registers[6][10] ),
    .A1(_3113_),
    .S(_3315_),
    .X(_3316_));
 sky130_fd_sc_hd__buf_1 _6801_ (.A(_3316_),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_2 _6802_ (.A0(\rf.registers[6][11] ),
    .A1(_3116_),
    .S(_3315_),
    .X(_3317_));
 sky130_fd_sc_hd__buf_1 _6803_ (.A(_3317_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_2 _6804_ (.A0(\rf.registers[6][12] ),
    .A1(_3118_),
    .S(_3315_),
    .X(_3318_));
 sky130_fd_sc_hd__buf_1 _6805_ (.A(_3318_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_2 _6806_ (.A0(\rf.registers[6][13] ),
    .A1(_3120_),
    .S(_3315_),
    .X(_3319_));
 sky130_fd_sc_hd__buf_1 _6807_ (.A(_3319_),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_2 _6808_ (.A0(\rf.registers[6][14] ),
    .A1(_3122_),
    .S(_3315_),
    .X(_3320_));
 sky130_fd_sc_hd__buf_1 _6809_ (.A(_3320_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_2 _6810_ (.A0(\rf.registers[6][15] ),
    .A1(_3124_),
    .S(_3315_),
    .X(_3321_));
 sky130_fd_sc_hd__buf_1 _6811_ (.A(_3321_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_2 _6812_ (.A0(\rf.registers[6][16] ),
    .A1(_3126_),
    .S(_3315_),
    .X(_3322_));
 sky130_fd_sc_hd__buf_1 _6813_ (.A(_3322_),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_2 _6814_ (.A0(\rf.registers[6][17] ),
    .A1(_3128_),
    .S(_3315_),
    .X(_3323_));
 sky130_fd_sc_hd__buf_1 _6815_ (.A(_3323_),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_2 _6816_ (.A0(\rf.registers[6][18] ),
    .A1(_3130_),
    .S(_3315_),
    .X(_3324_));
 sky130_fd_sc_hd__buf_1 _6817_ (.A(_3324_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_2 _6818_ (.A0(\rf.registers[6][19] ),
    .A1(_3132_),
    .S(_3315_),
    .X(_3325_));
 sky130_fd_sc_hd__buf_1 _6819_ (.A(_3325_),
    .X(_0969_));
 sky130_fd_sc_hd__buf_1 _6820_ (.A(_3303_),
    .X(_3326_));
 sky130_fd_sc_hd__mux2_2 _6821_ (.A0(\rf.registers[6][20] ),
    .A1(_3134_),
    .S(_3326_),
    .X(_3327_));
 sky130_fd_sc_hd__buf_1 _6822_ (.A(_3327_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_2 _6823_ (.A0(\rf.registers[6][21] ),
    .A1(_3137_),
    .S(_3326_),
    .X(_3328_));
 sky130_fd_sc_hd__buf_1 _6824_ (.A(_3328_),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_2 _6825_ (.A0(\rf.registers[6][22] ),
    .A1(_3139_),
    .S(_3326_),
    .X(_3329_));
 sky130_fd_sc_hd__buf_1 _6826_ (.A(_3329_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_2 _6827_ (.A0(\rf.registers[6][23] ),
    .A1(_3141_),
    .S(_3326_),
    .X(_3330_));
 sky130_fd_sc_hd__buf_1 _6828_ (.A(_3330_),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_2 _6829_ (.A0(\rf.registers[6][24] ),
    .A1(_3143_),
    .S(_3326_),
    .X(_3331_));
 sky130_fd_sc_hd__buf_1 _6830_ (.A(_3331_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_2 _6831_ (.A0(\rf.registers[6][25] ),
    .A1(_3145_),
    .S(_3326_),
    .X(_3332_));
 sky130_fd_sc_hd__buf_1 _6832_ (.A(_3332_),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_2 _6833_ (.A0(\rf.registers[6][26] ),
    .A1(_3002_),
    .S(_3326_),
    .X(_3333_));
 sky130_fd_sc_hd__buf_1 _6834_ (.A(_3333_),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_2 _6835_ (.A0(\rf.registers[6][27] ),
    .A1(_3009_),
    .S(_3326_),
    .X(_3334_));
 sky130_fd_sc_hd__buf_1 _6836_ (.A(_3334_),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_2 _6837_ (.A0(\rf.registers[6][28] ),
    .A1(_3011_),
    .S(_3326_),
    .X(_3335_));
 sky130_fd_sc_hd__buf_1 _6838_ (.A(_3335_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_2 _6839_ (.A0(\rf.registers[6][29] ),
    .A1(_3013_),
    .S(_3326_),
    .X(_3336_));
 sky130_fd_sc_hd__buf_1 _6840_ (.A(_3336_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_2 _6841_ (.A0(\rf.registers[6][30] ),
    .A1(_3015_),
    .S(_3303_),
    .X(_3337_));
 sky130_fd_sc_hd__buf_1 _6842_ (.A(_3337_),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_2 _6843_ (.A0(\rf.registers[6][31] ),
    .A1(_3017_),
    .S(_3303_),
    .X(_3338_));
 sky130_fd_sc_hd__buf_1 _6844_ (.A(_3338_),
    .X(_0981_));
 sky130_fd_sc_hd__nor2_2 _6845_ (.A(_3091_),
    .B(_3302_),
    .Y(_3339_));
 sky130_fd_sc_hd__buf_1 _6846_ (.A(_3339_),
    .X(_3340_));
 sky130_fd_sc_hd__mux2_2 _6847_ (.A0(\rf.registers[5][0] ),
    .A1(_3089_),
    .S(_3340_),
    .X(_3341_));
 sky130_fd_sc_hd__buf_1 _6848_ (.A(_3341_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_2 _6849_ (.A0(\rf.registers[5][1] ),
    .A1(_3095_),
    .S(_3340_),
    .X(_3342_));
 sky130_fd_sc_hd__buf_1 _6850_ (.A(_3342_),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_2 _6851_ (.A0(\rf.registers[5][2] ),
    .A1(_3097_),
    .S(_3340_),
    .X(_3343_));
 sky130_fd_sc_hd__buf_1 _6852_ (.A(_3343_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_2 _6853_ (.A0(\rf.registers[5][3] ),
    .A1(_3099_),
    .S(_3340_),
    .X(_3344_));
 sky130_fd_sc_hd__buf_1 _6854_ (.A(_3344_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_2 _6855_ (.A0(\rf.registers[5][4] ),
    .A1(_3101_),
    .S(_3340_),
    .X(_3345_));
 sky130_fd_sc_hd__buf_1 _6856_ (.A(_3345_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_2 _6857_ (.A0(\rf.registers[5][5] ),
    .A1(_3103_),
    .S(_3340_),
    .X(_3346_));
 sky130_fd_sc_hd__buf_1 _6858_ (.A(_3346_),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_2 _6859_ (.A0(\rf.registers[5][6] ),
    .A1(_3105_),
    .S(_3340_),
    .X(_3347_));
 sky130_fd_sc_hd__buf_1 _6860_ (.A(_3347_),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_2 _6861_ (.A0(\rf.registers[5][7] ),
    .A1(_3107_),
    .S(_3340_),
    .X(_3348_));
 sky130_fd_sc_hd__buf_1 _6862_ (.A(_3348_),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_2 _6863_ (.A0(\rf.registers[5][8] ),
    .A1(_3109_),
    .S(_3340_),
    .X(_3349_));
 sky130_fd_sc_hd__buf_1 _6864_ (.A(_3349_),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_2 _6865_ (.A0(\rf.registers[5][9] ),
    .A1(_3111_),
    .S(_3340_),
    .X(_3350_));
 sky130_fd_sc_hd__buf_1 _6866_ (.A(_3350_),
    .X(_0991_));
 sky130_fd_sc_hd__buf_1 _6867_ (.A(_3339_),
    .X(_3351_));
 sky130_fd_sc_hd__mux2_2 _6868_ (.A0(\rf.registers[5][10] ),
    .A1(_3113_),
    .S(_3351_),
    .X(_3352_));
 sky130_fd_sc_hd__buf_1 _6869_ (.A(_3352_),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_2 _6870_ (.A0(\rf.registers[5][11] ),
    .A1(_3116_),
    .S(_3351_),
    .X(_3353_));
 sky130_fd_sc_hd__buf_1 _6871_ (.A(_3353_),
    .X(_0993_));
 sky130_fd_sc_hd__mux2_2 _6872_ (.A0(\rf.registers[5][12] ),
    .A1(_3118_),
    .S(_3351_),
    .X(_3354_));
 sky130_fd_sc_hd__buf_1 _6873_ (.A(_3354_),
    .X(_0994_));
 sky130_fd_sc_hd__mux2_2 _6874_ (.A0(\rf.registers[5][13] ),
    .A1(_3120_),
    .S(_3351_),
    .X(_3355_));
 sky130_fd_sc_hd__buf_1 _6875_ (.A(_3355_),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_2 _6876_ (.A0(\rf.registers[5][14] ),
    .A1(_3122_),
    .S(_3351_),
    .X(_3356_));
 sky130_fd_sc_hd__buf_1 _6877_ (.A(_3356_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_2 _6878_ (.A0(\rf.registers[5][15] ),
    .A1(_3124_),
    .S(_3351_),
    .X(_3357_));
 sky130_fd_sc_hd__buf_1 _6879_ (.A(_3357_),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_2 _6880_ (.A0(\rf.registers[5][16] ),
    .A1(_3126_),
    .S(_3351_),
    .X(_3358_));
 sky130_fd_sc_hd__buf_1 _6881_ (.A(_3358_),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_2 _6882_ (.A0(\rf.registers[5][17] ),
    .A1(_3128_),
    .S(_3351_),
    .X(_3359_));
 sky130_fd_sc_hd__buf_1 _6883_ (.A(_3359_),
    .X(_0999_));
 sky130_fd_sc_hd__mux2_2 _6884_ (.A0(\rf.registers[5][18] ),
    .A1(_3130_),
    .S(_3351_),
    .X(_3360_));
 sky130_fd_sc_hd__buf_1 _6885_ (.A(_3360_),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_2 _6886_ (.A0(\rf.registers[5][19] ),
    .A1(_3132_),
    .S(_3351_),
    .X(_3361_));
 sky130_fd_sc_hd__buf_1 _6887_ (.A(_3361_),
    .X(_1001_));
 sky130_fd_sc_hd__buf_1 _6888_ (.A(_3339_),
    .X(_3362_));
 sky130_fd_sc_hd__mux2_2 _6889_ (.A0(\rf.registers[5][20] ),
    .A1(_3134_),
    .S(_3362_),
    .X(_3363_));
 sky130_fd_sc_hd__buf_1 _6890_ (.A(_3363_),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_2 _6891_ (.A0(\rf.registers[5][21] ),
    .A1(_3137_),
    .S(_3362_),
    .X(_3364_));
 sky130_fd_sc_hd__buf_1 _6892_ (.A(_3364_),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_2 _6893_ (.A0(\rf.registers[5][22] ),
    .A1(_3139_),
    .S(_3362_),
    .X(_3365_));
 sky130_fd_sc_hd__buf_1 _6894_ (.A(_3365_),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_2 _6895_ (.A0(\rf.registers[5][23] ),
    .A1(_3141_),
    .S(_3362_),
    .X(_3366_));
 sky130_fd_sc_hd__buf_1 _6896_ (.A(_3366_),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_2 _6897_ (.A0(\rf.registers[5][24] ),
    .A1(_3143_),
    .S(_3362_),
    .X(_3367_));
 sky130_fd_sc_hd__buf_1 _6898_ (.A(_3367_),
    .X(_1006_));
 sky130_fd_sc_hd__mux2_2 _6899_ (.A0(\rf.registers[5][25] ),
    .A1(_3145_),
    .S(_3362_),
    .X(_3368_));
 sky130_fd_sc_hd__buf_1 _6900_ (.A(_3368_),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_2 _6901_ (.A0(\rf.registers[5][26] ),
    .A1(_3002_),
    .S(_3362_),
    .X(_3369_));
 sky130_fd_sc_hd__buf_1 _6902_ (.A(_3369_),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_2 _6903_ (.A0(\rf.registers[5][27] ),
    .A1(_3009_),
    .S(_3362_),
    .X(_3370_));
 sky130_fd_sc_hd__buf_1 _6904_ (.A(_3370_),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_2 _6905_ (.A0(\rf.registers[5][28] ),
    .A1(_3011_),
    .S(_3362_),
    .X(_3371_));
 sky130_fd_sc_hd__buf_1 _6906_ (.A(_3371_),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_2 _6907_ (.A0(\rf.registers[5][29] ),
    .A1(_3013_),
    .S(_3362_),
    .X(_3372_));
 sky130_fd_sc_hd__buf_1 _6908_ (.A(_3372_),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_2 _6909_ (.A0(\rf.registers[5][30] ),
    .A1(_3015_),
    .S(_3339_),
    .X(_3373_));
 sky130_fd_sc_hd__buf_1 _6910_ (.A(_3373_),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_2 _6911_ (.A0(\rf.registers[5][31] ),
    .A1(_3017_),
    .S(_3339_),
    .X(_3374_));
 sky130_fd_sc_hd__buf_1 _6912_ (.A(_3374_),
    .X(_1013_));
 sky130_fd_sc_hd__nor2_2 _6913_ (.A(_3155_),
    .B(_3302_),
    .Y(_3375_));
 sky130_fd_sc_hd__buf_1 _6914_ (.A(_3375_),
    .X(_3376_));
 sky130_fd_sc_hd__mux2_2 _6915_ (.A0(\rf.registers[4][0] ),
    .A1(_3089_),
    .S(_3376_),
    .X(_3377_));
 sky130_fd_sc_hd__buf_1 _6916_ (.A(_3377_),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_2 _6917_ (.A0(\rf.registers[4][1] ),
    .A1(_3095_),
    .S(_3376_),
    .X(_3378_));
 sky130_fd_sc_hd__buf_1 _6918_ (.A(_3378_),
    .X(_1015_));
 sky130_fd_sc_hd__mux2_2 _6919_ (.A0(\rf.registers[4][2] ),
    .A1(_3097_),
    .S(_3376_),
    .X(_3379_));
 sky130_fd_sc_hd__buf_1 _6920_ (.A(_3379_),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_2 _6921_ (.A0(\rf.registers[4][3] ),
    .A1(_3099_),
    .S(_3376_),
    .X(_3380_));
 sky130_fd_sc_hd__buf_1 _6922_ (.A(_3380_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_2 _6923_ (.A0(\rf.registers[4][4] ),
    .A1(_3101_),
    .S(_3376_),
    .X(_3381_));
 sky130_fd_sc_hd__buf_1 _6924_ (.A(_3381_),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_2 _6925_ (.A0(\rf.registers[4][5] ),
    .A1(_3103_),
    .S(_3376_),
    .X(_3382_));
 sky130_fd_sc_hd__buf_1 _6926_ (.A(_3382_),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_2 _6927_ (.A0(\rf.registers[4][6] ),
    .A1(_3105_),
    .S(_3376_),
    .X(_3383_));
 sky130_fd_sc_hd__buf_1 _6928_ (.A(_3383_),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_2 _6929_ (.A0(\rf.registers[4][7] ),
    .A1(_3107_),
    .S(_3376_),
    .X(_3384_));
 sky130_fd_sc_hd__buf_1 _6930_ (.A(_3384_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_2 _6931_ (.A0(\rf.registers[4][8] ),
    .A1(_3109_),
    .S(_3376_),
    .X(_3385_));
 sky130_fd_sc_hd__buf_1 _6932_ (.A(_3385_),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_2 _6933_ (.A0(\rf.registers[4][9] ),
    .A1(_3111_),
    .S(_3376_),
    .X(_3386_));
 sky130_fd_sc_hd__buf_1 _6934_ (.A(_3386_),
    .X(_1023_));
 sky130_fd_sc_hd__buf_1 _6935_ (.A(_3375_),
    .X(_3387_));
 sky130_fd_sc_hd__mux2_2 _6936_ (.A0(\rf.registers[4][10] ),
    .A1(_3113_),
    .S(_3387_),
    .X(_3388_));
 sky130_fd_sc_hd__buf_1 _6937_ (.A(_3388_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_2 _6938_ (.A0(\rf.registers[4][11] ),
    .A1(_3116_),
    .S(_3387_),
    .X(_3389_));
 sky130_fd_sc_hd__buf_1 _6939_ (.A(_3389_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_2 _6940_ (.A0(\rf.registers[4][12] ),
    .A1(_3118_),
    .S(_3387_),
    .X(_3390_));
 sky130_fd_sc_hd__buf_1 _6941_ (.A(_3390_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_2 _6942_ (.A0(\rf.registers[4][13] ),
    .A1(_3120_),
    .S(_3387_),
    .X(_3391_));
 sky130_fd_sc_hd__buf_1 _6943_ (.A(_3391_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_2 _6944_ (.A0(\rf.registers[4][14] ),
    .A1(_3122_),
    .S(_3387_),
    .X(_3392_));
 sky130_fd_sc_hd__buf_1 _6945_ (.A(_3392_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_2 _6946_ (.A0(\rf.registers[4][15] ),
    .A1(_3124_),
    .S(_3387_),
    .X(_3393_));
 sky130_fd_sc_hd__buf_1 _6947_ (.A(_3393_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_2 _6948_ (.A0(\rf.registers[4][16] ),
    .A1(_3126_),
    .S(_3387_),
    .X(_3394_));
 sky130_fd_sc_hd__buf_1 _6949_ (.A(_3394_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_2 _6950_ (.A0(\rf.registers[4][17] ),
    .A1(_3128_),
    .S(_3387_),
    .X(_3395_));
 sky130_fd_sc_hd__buf_1 _6951_ (.A(_3395_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_2 _6952_ (.A0(\rf.registers[4][18] ),
    .A1(_3130_),
    .S(_3387_),
    .X(_3396_));
 sky130_fd_sc_hd__buf_1 _6953_ (.A(_3396_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_2 _6954_ (.A0(\rf.registers[4][19] ),
    .A1(_3132_),
    .S(_3387_),
    .X(_3397_));
 sky130_fd_sc_hd__buf_1 _6955_ (.A(_3397_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_1 _6956_ (.A(_3375_),
    .X(_3398_));
 sky130_fd_sc_hd__mux2_2 _6957_ (.A0(\rf.registers[4][20] ),
    .A1(_3134_),
    .S(_3398_),
    .X(_3399_));
 sky130_fd_sc_hd__buf_1 _6958_ (.A(_3399_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_2 _6959_ (.A0(\rf.registers[4][21] ),
    .A1(_3137_),
    .S(_3398_),
    .X(_3400_));
 sky130_fd_sc_hd__buf_1 _6960_ (.A(_3400_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_2 _6961_ (.A0(\rf.registers[4][22] ),
    .A1(_3139_),
    .S(_3398_),
    .X(_3401_));
 sky130_fd_sc_hd__buf_1 _6962_ (.A(_3401_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_2 _6963_ (.A0(\rf.registers[4][23] ),
    .A1(_3141_),
    .S(_3398_),
    .X(_3402_));
 sky130_fd_sc_hd__buf_1 _6964_ (.A(_3402_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_2 _6965_ (.A0(\rf.registers[4][24] ),
    .A1(_3143_),
    .S(_3398_),
    .X(_3403_));
 sky130_fd_sc_hd__buf_1 _6966_ (.A(_3403_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_2 _6967_ (.A0(\rf.registers[4][25] ),
    .A1(_3145_),
    .S(_3398_),
    .X(_3404_));
 sky130_fd_sc_hd__buf_1 _6968_ (.A(_3404_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_2 _6969_ (.A0(\rf.registers[4][26] ),
    .A1(_3002_),
    .S(_3398_),
    .X(_3405_));
 sky130_fd_sc_hd__buf_1 _6970_ (.A(_3405_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_2 _6971_ (.A0(\rf.registers[4][27] ),
    .A1(_3009_),
    .S(_3398_),
    .X(_3406_));
 sky130_fd_sc_hd__buf_1 _6972_ (.A(_3406_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_2 _6973_ (.A0(\rf.registers[4][28] ),
    .A1(_3011_),
    .S(_3398_),
    .X(_3407_));
 sky130_fd_sc_hd__buf_1 _6974_ (.A(_3407_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_2 _6975_ (.A0(\rf.registers[4][29] ),
    .A1(_3013_),
    .S(_3398_),
    .X(_3408_));
 sky130_fd_sc_hd__buf_1 _6976_ (.A(_3408_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_2 _6977_ (.A0(\rf.registers[4][30] ),
    .A1(_3015_),
    .S(_3375_),
    .X(_3409_));
 sky130_fd_sc_hd__buf_1 _6978_ (.A(_3409_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_2 _6979_ (.A0(\rf.registers[4][31] ),
    .A1(_3017_),
    .S(_3375_),
    .X(_3410_));
 sky130_fd_sc_hd__buf_1 _6980_ (.A(_3410_),
    .X(_0021_));
 sky130_fd_sc_hd__nand3_2 _6981_ (.A(A3[1]),
    .B(A3[0]),
    .C(WE3),
    .Y(_3411_));
 sky130_fd_sc_hd__nor2_2 _6982_ (.A(_3090_),
    .B(_3411_),
    .Y(_3412_));
 sky130_fd_sc_hd__buf_1 _6983_ (.A(_3412_),
    .X(_3413_));
 sky130_fd_sc_hd__mux2_2 _6984_ (.A0(\rf.registers[19][0] ),
    .A1(_3089_),
    .S(_3413_),
    .X(_3414_));
 sky130_fd_sc_hd__buf_1 _6985_ (.A(_3414_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_2 _6986_ (.A0(\rf.registers[19][1] ),
    .A1(_3095_),
    .S(_3413_),
    .X(_3415_));
 sky130_fd_sc_hd__buf_1 _6987_ (.A(_3415_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_2 _6988_ (.A0(\rf.registers[19][2] ),
    .A1(_3097_),
    .S(_3413_),
    .X(_3416_));
 sky130_fd_sc_hd__buf_1 _6989_ (.A(_3416_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_2 _6990_ (.A0(\rf.registers[19][3] ),
    .A1(_3099_),
    .S(_3413_),
    .X(_3417_));
 sky130_fd_sc_hd__buf_1 _6991_ (.A(_3417_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_2 _6992_ (.A0(\rf.registers[19][4] ),
    .A1(_3101_),
    .S(_3413_),
    .X(_3418_));
 sky130_fd_sc_hd__buf_1 _6993_ (.A(_3418_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_2 _6994_ (.A0(\rf.registers[19][5] ),
    .A1(_3103_),
    .S(_3413_),
    .X(_3419_));
 sky130_fd_sc_hd__buf_1 _6995_ (.A(_3419_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_2 _6996_ (.A0(\rf.registers[19][6] ),
    .A1(_3105_),
    .S(_3413_),
    .X(_3420_));
 sky130_fd_sc_hd__buf_1 _6997_ (.A(_3420_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_2 _6998_ (.A0(\rf.registers[19][7] ),
    .A1(_3107_),
    .S(_3413_),
    .X(_3421_));
 sky130_fd_sc_hd__buf_1 _6999_ (.A(_3421_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_2 _7000_ (.A0(\rf.registers[19][8] ),
    .A1(_3109_),
    .S(_3413_),
    .X(_3422_));
 sky130_fd_sc_hd__buf_1 _7001_ (.A(_3422_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_2 _7002_ (.A0(\rf.registers[19][9] ),
    .A1(_3111_),
    .S(_3413_),
    .X(_3423_));
 sky130_fd_sc_hd__buf_1 _7003_ (.A(_3423_),
    .X(_0031_));
 sky130_fd_sc_hd__buf_1 _7004_ (.A(_3412_),
    .X(_3424_));
 sky130_fd_sc_hd__mux2_2 _7005_ (.A0(\rf.registers[19][10] ),
    .A1(_3113_),
    .S(_3424_),
    .X(_3425_));
 sky130_fd_sc_hd__buf_1 _7006_ (.A(_3425_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_2 _7007_ (.A0(\rf.registers[19][11] ),
    .A1(_3116_),
    .S(_3424_),
    .X(_3426_));
 sky130_fd_sc_hd__buf_1 _7008_ (.A(_3426_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_2 _7009_ (.A0(\rf.registers[19][12] ),
    .A1(_3118_),
    .S(_3424_),
    .X(_3427_));
 sky130_fd_sc_hd__buf_1 _7010_ (.A(_3427_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_2 _7011_ (.A0(\rf.registers[19][13] ),
    .A1(_3120_),
    .S(_3424_),
    .X(_3428_));
 sky130_fd_sc_hd__buf_1 _7012_ (.A(_3428_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_2 _7013_ (.A0(\rf.registers[19][14] ),
    .A1(_3122_),
    .S(_3424_),
    .X(_3429_));
 sky130_fd_sc_hd__buf_1 _7014_ (.A(_3429_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_2 _7015_ (.A0(\rf.registers[19][15] ),
    .A1(_3124_),
    .S(_3424_),
    .X(_3430_));
 sky130_fd_sc_hd__buf_1 _7016_ (.A(_3430_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_2 _7017_ (.A0(\rf.registers[19][16] ),
    .A1(_3126_),
    .S(_3424_),
    .X(_3431_));
 sky130_fd_sc_hd__buf_1 _7018_ (.A(_3431_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_2 _7019_ (.A0(\rf.registers[19][17] ),
    .A1(_3128_),
    .S(_3424_),
    .X(_3432_));
 sky130_fd_sc_hd__buf_1 _7020_ (.A(_3432_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_2 _7021_ (.A0(\rf.registers[19][18] ),
    .A1(_3130_),
    .S(_3424_),
    .X(_3433_));
 sky130_fd_sc_hd__buf_1 _7022_ (.A(_3433_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_2 _7023_ (.A0(\rf.registers[19][19] ),
    .A1(_3132_),
    .S(_3424_),
    .X(_3434_));
 sky130_fd_sc_hd__buf_1 _7024_ (.A(_3434_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_1 _7025_ (.A(_3412_),
    .X(_3435_));
 sky130_fd_sc_hd__mux2_2 _7026_ (.A0(\rf.registers[19][20] ),
    .A1(_3134_),
    .S(_3435_),
    .X(_3436_));
 sky130_fd_sc_hd__buf_1 _7027_ (.A(_3436_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_2 _7028_ (.A0(\rf.registers[19][21] ),
    .A1(_3137_),
    .S(_3435_),
    .X(_3437_));
 sky130_fd_sc_hd__buf_1 _7029_ (.A(_3437_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_2 _7030_ (.A0(\rf.registers[19][22] ),
    .A1(_3139_),
    .S(_3435_),
    .X(_3438_));
 sky130_fd_sc_hd__buf_1 _7031_ (.A(_3438_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_2 _7032_ (.A0(\rf.registers[19][23] ),
    .A1(_3141_),
    .S(_3435_),
    .X(_3439_));
 sky130_fd_sc_hd__buf_1 _7033_ (.A(_3439_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_2 _7034_ (.A0(\rf.registers[19][24] ),
    .A1(_3143_),
    .S(_3435_),
    .X(_3440_));
 sky130_fd_sc_hd__buf_1 _7035_ (.A(_3440_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_2 _7036_ (.A0(\rf.registers[19][25] ),
    .A1(_3145_),
    .S(_3435_),
    .X(_3441_));
 sky130_fd_sc_hd__buf_1 _7037_ (.A(_3441_),
    .X(_0047_));
 sky130_fd_sc_hd__buf_1 _7038_ (.A(WD3[26]),
    .X(_3442_));
 sky130_fd_sc_hd__mux2_2 _7039_ (.A0(\rf.registers[19][26] ),
    .A1(_3442_),
    .S(_3435_),
    .X(_3443_));
 sky130_fd_sc_hd__buf_1 _7040_ (.A(_3443_),
    .X(_0048_));
 sky130_fd_sc_hd__buf_1 _7041_ (.A(WD3[27]),
    .X(_3444_));
 sky130_fd_sc_hd__mux2_2 _7042_ (.A0(\rf.registers[19][27] ),
    .A1(_3444_),
    .S(_3435_),
    .X(_3445_));
 sky130_fd_sc_hd__buf_1 _7043_ (.A(_3445_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_1 _7044_ (.A(WD3[28]),
    .X(_3446_));
 sky130_fd_sc_hd__mux2_2 _7045_ (.A0(\rf.registers[19][28] ),
    .A1(_3446_),
    .S(_3435_),
    .X(_3447_));
 sky130_fd_sc_hd__buf_1 _7046_ (.A(_3447_),
    .X(_0050_));
 sky130_fd_sc_hd__buf_1 _7047_ (.A(WD3[29]),
    .X(_3448_));
 sky130_fd_sc_hd__mux2_2 _7048_ (.A0(\rf.registers[19][29] ),
    .A1(_3448_),
    .S(_3435_),
    .X(_3449_));
 sky130_fd_sc_hd__buf_1 _7049_ (.A(_3449_),
    .X(_0051_));
 sky130_fd_sc_hd__buf_1 _7050_ (.A(WD3[30]),
    .X(_3450_));
 sky130_fd_sc_hd__mux2_2 _7051_ (.A0(\rf.registers[19][30] ),
    .A1(_3450_),
    .S(_3412_),
    .X(_3451_));
 sky130_fd_sc_hd__buf_1 _7052_ (.A(_3451_),
    .X(_0052_));
 sky130_fd_sc_hd__buf_1 _7053_ (.A(WD3[31]),
    .X(_3452_));
 sky130_fd_sc_hd__mux2_2 _7054_ (.A0(\rf.registers[19][31] ),
    .A1(_3452_),
    .S(_3412_),
    .X(_3453_));
 sky130_fd_sc_hd__buf_1 _7055_ (.A(_3453_),
    .X(_0053_));
 sky130_fd_sc_hd__buf_1 _7056_ (.A(WD3[0]),
    .X(_3454_));
 sky130_fd_sc_hd__nor2_2 _7057_ (.A(_3153_),
    .B(_3411_),
    .Y(_3455_));
 sky130_fd_sc_hd__buf_1 _7058_ (.A(_3455_),
    .X(_3456_));
 sky130_fd_sc_hd__mux2_2 _7059_ (.A0(\rf.registers[3][0] ),
    .A1(_3454_),
    .S(_3456_),
    .X(_3457_));
 sky130_fd_sc_hd__buf_1 _7060_ (.A(_3457_),
    .X(_0054_));
 sky130_fd_sc_hd__buf_1 _7061_ (.A(WD3[1]),
    .X(_3458_));
 sky130_fd_sc_hd__mux2_2 _7062_ (.A0(\rf.registers[3][1] ),
    .A1(_3458_),
    .S(_3456_),
    .X(_3459_));
 sky130_fd_sc_hd__buf_1 _7063_ (.A(_3459_),
    .X(_0055_));
 sky130_fd_sc_hd__buf_1 _7064_ (.A(WD3[2]),
    .X(_3460_));
 sky130_fd_sc_hd__mux2_2 _7065_ (.A0(\rf.registers[3][2] ),
    .A1(_3460_),
    .S(_3456_),
    .X(_3461_));
 sky130_fd_sc_hd__buf_1 _7066_ (.A(_3461_),
    .X(_0056_));
 sky130_fd_sc_hd__buf_1 _7067_ (.A(WD3[3]),
    .X(_3462_));
 sky130_fd_sc_hd__mux2_2 _7068_ (.A0(\rf.registers[3][3] ),
    .A1(_3462_),
    .S(_3456_),
    .X(_3463_));
 sky130_fd_sc_hd__buf_1 _7069_ (.A(_3463_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_1 _7070_ (.A(WD3[4]),
    .X(_3464_));
 sky130_fd_sc_hd__mux2_2 _7071_ (.A0(\rf.registers[3][4] ),
    .A1(_3464_),
    .S(_3456_),
    .X(_3465_));
 sky130_fd_sc_hd__buf_1 _7072_ (.A(_3465_),
    .X(_0058_));
 sky130_fd_sc_hd__buf_1 _7073_ (.A(WD3[5]),
    .X(_3466_));
 sky130_fd_sc_hd__mux2_2 _7074_ (.A0(\rf.registers[3][5] ),
    .A1(_3466_),
    .S(_3456_),
    .X(_3467_));
 sky130_fd_sc_hd__buf_1 _7075_ (.A(_3467_),
    .X(_0059_));
 sky130_fd_sc_hd__buf_1 _7076_ (.A(WD3[6]),
    .X(_3468_));
 sky130_fd_sc_hd__mux2_2 _7077_ (.A0(\rf.registers[3][6] ),
    .A1(_3468_),
    .S(_3456_),
    .X(_3469_));
 sky130_fd_sc_hd__buf_1 _7078_ (.A(_3469_),
    .X(_0060_));
 sky130_fd_sc_hd__buf_1 _7079_ (.A(WD3[7]),
    .X(_3470_));
 sky130_fd_sc_hd__mux2_2 _7080_ (.A0(\rf.registers[3][7] ),
    .A1(_3470_),
    .S(_3456_),
    .X(_3471_));
 sky130_fd_sc_hd__buf_1 _7081_ (.A(_3471_),
    .X(_0061_));
 sky130_fd_sc_hd__buf_1 _7082_ (.A(WD3[8]),
    .X(_3472_));
 sky130_fd_sc_hd__mux2_2 _7083_ (.A0(\rf.registers[3][8] ),
    .A1(_3472_),
    .S(_3456_),
    .X(_3473_));
 sky130_fd_sc_hd__buf_1 _7084_ (.A(_3473_),
    .X(_0062_));
 sky130_fd_sc_hd__buf_1 _7085_ (.A(WD3[9]),
    .X(_3474_));
 sky130_fd_sc_hd__mux2_2 _7086_ (.A0(\rf.registers[3][9] ),
    .A1(_3474_),
    .S(_3456_),
    .X(_3475_));
 sky130_fd_sc_hd__buf_1 _7087_ (.A(_3475_),
    .X(_0063_));
 sky130_fd_sc_hd__buf_1 _7088_ (.A(WD3[10]),
    .X(_3476_));
 sky130_fd_sc_hd__buf_1 _7089_ (.A(_3455_),
    .X(_3477_));
 sky130_fd_sc_hd__mux2_2 _7090_ (.A0(\rf.registers[3][10] ),
    .A1(_3476_),
    .S(_3477_),
    .X(_3478_));
 sky130_fd_sc_hd__buf_1 _7091_ (.A(_3478_),
    .X(_0064_));
 sky130_fd_sc_hd__buf_1 _7092_ (.A(WD3[11]),
    .X(_3479_));
 sky130_fd_sc_hd__mux2_2 _7093_ (.A0(\rf.registers[3][11] ),
    .A1(_3479_),
    .S(_3477_),
    .X(_3480_));
 sky130_fd_sc_hd__buf_1 _7094_ (.A(_3480_),
    .X(_0065_));
 sky130_fd_sc_hd__buf_1 _7095_ (.A(WD3[12]),
    .X(_3481_));
 sky130_fd_sc_hd__mux2_2 _7096_ (.A0(\rf.registers[3][12] ),
    .A1(_3481_),
    .S(_3477_),
    .X(_3482_));
 sky130_fd_sc_hd__buf_1 _7097_ (.A(_3482_),
    .X(_0066_));
 sky130_fd_sc_hd__buf_1 _7098_ (.A(WD3[13]),
    .X(_3483_));
 sky130_fd_sc_hd__mux2_2 _7099_ (.A0(\rf.registers[3][13] ),
    .A1(_3483_),
    .S(_3477_),
    .X(_3484_));
 sky130_fd_sc_hd__buf_1 _7100_ (.A(_3484_),
    .X(_0067_));
 sky130_fd_sc_hd__buf_1 _7101_ (.A(WD3[14]),
    .X(_3485_));
 sky130_fd_sc_hd__mux2_2 _7102_ (.A0(\rf.registers[3][14] ),
    .A1(_3485_),
    .S(_3477_),
    .X(_3486_));
 sky130_fd_sc_hd__buf_1 _7103_ (.A(_3486_),
    .X(_0068_));
 sky130_fd_sc_hd__buf_1 _7104_ (.A(WD3[15]),
    .X(_3487_));
 sky130_fd_sc_hd__mux2_2 _7105_ (.A0(\rf.registers[3][15] ),
    .A1(_3487_),
    .S(_3477_),
    .X(_3488_));
 sky130_fd_sc_hd__buf_1 _7106_ (.A(_3488_),
    .X(_0069_));
 sky130_fd_sc_hd__buf_1 _7107_ (.A(WD3[16]),
    .X(_3489_));
 sky130_fd_sc_hd__mux2_2 _7108_ (.A0(\rf.registers[3][16] ),
    .A1(_3489_),
    .S(_3477_),
    .X(_3490_));
 sky130_fd_sc_hd__buf_1 _7109_ (.A(_3490_),
    .X(_0070_));
 sky130_fd_sc_hd__buf_1 _7110_ (.A(WD3[17]),
    .X(_3491_));
 sky130_fd_sc_hd__mux2_2 _7111_ (.A0(\rf.registers[3][17] ),
    .A1(_3491_),
    .S(_3477_),
    .X(_3492_));
 sky130_fd_sc_hd__buf_1 _7112_ (.A(_3492_),
    .X(_0071_));
 sky130_fd_sc_hd__buf_1 _7113_ (.A(WD3[18]),
    .X(_3493_));
 sky130_fd_sc_hd__mux2_2 _7114_ (.A0(\rf.registers[3][18] ),
    .A1(_3493_),
    .S(_3477_),
    .X(_3494_));
 sky130_fd_sc_hd__buf_1 _7115_ (.A(_3494_),
    .X(_0072_));
 sky130_fd_sc_hd__buf_1 _7116_ (.A(WD3[19]),
    .X(_3495_));
 sky130_fd_sc_hd__mux2_2 _7117_ (.A0(\rf.registers[3][19] ),
    .A1(_3495_),
    .S(_3477_),
    .X(_3496_));
 sky130_fd_sc_hd__buf_1 _7118_ (.A(_3496_),
    .X(_0073_));
 sky130_fd_sc_hd__buf_1 _7119_ (.A(WD3[20]),
    .X(_3497_));
 sky130_fd_sc_hd__buf_1 _7120_ (.A(_3455_),
    .X(_3498_));
 sky130_fd_sc_hd__mux2_2 _7121_ (.A0(\rf.registers[3][20] ),
    .A1(_3497_),
    .S(_3498_),
    .X(_3499_));
 sky130_fd_sc_hd__buf_1 _7122_ (.A(_3499_),
    .X(_0074_));
 sky130_fd_sc_hd__buf_1 _7123_ (.A(WD3[21]),
    .X(_3500_));
 sky130_fd_sc_hd__mux2_2 _7124_ (.A0(\rf.registers[3][21] ),
    .A1(_3500_),
    .S(_3498_),
    .X(_3501_));
 sky130_fd_sc_hd__buf_1 _7125_ (.A(_3501_),
    .X(_0075_));
 sky130_fd_sc_hd__buf_1 _7126_ (.A(WD3[22]),
    .X(_3502_));
 sky130_fd_sc_hd__mux2_2 _7127_ (.A0(\rf.registers[3][22] ),
    .A1(_3502_),
    .S(_3498_),
    .X(_3503_));
 sky130_fd_sc_hd__buf_1 _7128_ (.A(_3503_),
    .X(_0076_));
 sky130_fd_sc_hd__buf_1 _7129_ (.A(WD3[23]),
    .X(_3504_));
 sky130_fd_sc_hd__mux2_2 _7130_ (.A0(\rf.registers[3][23] ),
    .A1(_3504_),
    .S(_3498_),
    .X(_3505_));
 sky130_fd_sc_hd__buf_1 _7131_ (.A(_3505_),
    .X(_0077_));
 sky130_fd_sc_hd__buf_1 _7132_ (.A(WD3[24]),
    .X(_3506_));
 sky130_fd_sc_hd__mux2_2 _7133_ (.A0(\rf.registers[3][24] ),
    .A1(_3506_),
    .S(_3498_),
    .X(_3507_));
 sky130_fd_sc_hd__buf_1 _7134_ (.A(_3507_),
    .X(_0078_));
 sky130_fd_sc_hd__buf_1 _7135_ (.A(WD3[25]),
    .X(_3508_));
 sky130_fd_sc_hd__mux2_2 _7136_ (.A0(\rf.registers[3][25] ),
    .A1(_3508_),
    .S(_3498_),
    .X(_3509_));
 sky130_fd_sc_hd__buf_1 _7137_ (.A(_3509_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_2 _7138_ (.A0(\rf.registers[3][26] ),
    .A1(_3442_),
    .S(_3498_),
    .X(_3510_));
 sky130_fd_sc_hd__buf_1 _7139_ (.A(_3510_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_2 _7140_ (.A0(\rf.registers[3][27] ),
    .A1(_3444_),
    .S(_3498_),
    .X(_3511_));
 sky130_fd_sc_hd__buf_1 _7141_ (.A(_3511_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_2 _7142_ (.A0(\rf.registers[3][28] ),
    .A1(_3446_),
    .S(_3498_),
    .X(_3512_));
 sky130_fd_sc_hd__buf_1 _7143_ (.A(_3512_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_2 _7144_ (.A0(\rf.registers[3][29] ),
    .A1(_3448_),
    .S(_3498_),
    .X(_3513_));
 sky130_fd_sc_hd__buf_1 _7145_ (.A(_3513_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_2 _7146_ (.A0(\rf.registers[3][30] ),
    .A1(_3450_),
    .S(_3455_),
    .X(_3514_));
 sky130_fd_sc_hd__buf_1 _7147_ (.A(_3514_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_2 _7148_ (.A0(\rf.registers[3][31] ),
    .A1(_3452_),
    .S(_3455_),
    .X(_3515_));
 sky130_fd_sc_hd__buf_1 _7149_ (.A(_3515_),
    .X(_0085_));
 sky130_fd_sc_hd__nor2_2 _7150_ (.A(_3411_),
    .B(_3302_),
    .Y(_3516_));
 sky130_fd_sc_hd__buf_1 _7151_ (.A(_3516_),
    .X(_3517_));
 sky130_fd_sc_hd__mux2_2 _7152_ (.A0(\rf.registers[7][0] ),
    .A1(_3454_),
    .S(_3517_),
    .X(_3518_));
 sky130_fd_sc_hd__buf_1 _7153_ (.A(_3518_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_2 _7154_ (.A0(\rf.registers[7][1] ),
    .A1(_3458_),
    .S(_3517_),
    .X(_3519_));
 sky130_fd_sc_hd__buf_1 _7155_ (.A(_3519_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_2 _7156_ (.A0(\rf.registers[7][2] ),
    .A1(_3460_),
    .S(_3517_),
    .X(_3520_));
 sky130_fd_sc_hd__buf_1 _7157_ (.A(_3520_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_2 _7158_ (.A0(\rf.registers[7][3] ),
    .A1(_3462_),
    .S(_3517_),
    .X(_3521_));
 sky130_fd_sc_hd__buf_1 _7159_ (.A(_3521_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_2 _7160_ (.A0(\rf.registers[7][4] ),
    .A1(_3464_),
    .S(_3517_),
    .X(_3522_));
 sky130_fd_sc_hd__buf_1 _7161_ (.A(_3522_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_2 _7162_ (.A0(\rf.registers[7][5] ),
    .A1(_3466_),
    .S(_3517_),
    .X(_3523_));
 sky130_fd_sc_hd__buf_1 _7163_ (.A(_3523_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_2 _7164_ (.A0(\rf.registers[7][6] ),
    .A1(_3468_),
    .S(_3517_),
    .X(_3524_));
 sky130_fd_sc_hd__buf_1 _7165_ (.A(_3524_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_2 _7166_ (.A0(\rf.registers[7][7] ),
    .A1(_3470_),
    .S(_3517_),
    .X(_3525_));
 sky130_fd_sc_hd__buf_1 _7167_ (.A(_3525_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_2 _7168_ (.A0(\rf.registers[7][8] ),
    .A1(_3472_),
    .S(_3517_),
    .X(_3526_));
 sky130_fd_sc_hd__buf_1 _7169_ (.A(_3526_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_2 _7170_ (.A0(\rf.registers[7][9] ),
    .A1(_3474_),
    .S(_3517_),
    .X(_3527_));
 sky130_fd_sc_hd__buf_1 _7171_ (.A(_3527_),
    .X(_0095_));
 sky130_fd_sc_hd__buf_1 _7172_ (.A(_3516_),
    .X(_3528_));
 sky130_fd_sc_hd__mux2_2 _7173_ (.A0(\rf.registers[7][10] ),
    .A1(_3476_),
    .S(_3528_),
    .X(_3529_));
 sky130_fd_sc_hd__buf_1 _7174_ (.A(_3529_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_2 _7175_ (.A0(\rf.registers[7][11] ),
    .A1(_3479_),
    .S(_3528_),
    .X(_3530_));
 sky130_fd_sc_hd__buf_1 _7176_ (.A(_3530_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_2 _7177_ (.A0(\rf.registers[7][12] ),
    .A1(_3481_),
    .S(_3528_),
    .X(_3531_));
 sky130_fd_sc_hd__buf_1 _7178_ (.A(_3531_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_2 _7179_ (.A0(\rf.registers[7][13] ),
    .A1(_3483_),
    .S(_3528_),
    .X(_3532_));
 sky130_fd_sc_hd__buf_1 _7180_ (.A(_3532_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_2 _7181_ (.A0(\rf.registers[7][14] ),
    .A1(_3485_),
    .S(_3528_),
    .X(_3533_));
 sky130_fd_sc_hd__buf_1 _7182_ (.A(_3533_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_2 _7183_ (.A0(\rf.registers[7][15] ),
    .A1(_3487_),
    .S(_3528_),
    .X(_3534_));
 sky130_fd_sc_hd__buf_1 _7184_ (.A(_3534_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_2 _7185_ (.A0(\rf.registers[7][16] ),
    .A1(_3489_),
    .S(_3528_),
    .X(_3535_));
 sky130_fd_sc_hd__buf_1 _7186_ (.A(_3535_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_2 _7187_ (.A0(\rf.registers[7][17] ),
    .A1(_3491_),
    .S(_3528_),
    .X(_3536_));
 sky130_fd_sc_hd__buf_1 _7188_ (.A(_3536_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_2 _7189_ (.A0(\rf.registers[7][18] ),
    .A1(_3493_),
    .S(_3528_),
    .X(_3537_));
 sky130_fd_sc_hd__buf_1 _7190_ (.A(_3537_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_2 _7191_ (.A0(\rf.registers[7][19] ),
    .A1(_3495_),
    .S(_3528_),
    .X(_3538_));
 sky130_fd_sc_hd__buf_1 _7192_ (.A(_3538_),
    .X(_0105_));
 sky130_fd_sc_hd__buf_1 _7193_ (.A(_3516_),
    .X(_3539_));
 sky130_fd_sc_hd__mux2_2 _7194_ (.A0(\rf.registers[7][20] ),
    .A1(_3497_),
    .S(_3539_),
    .X(_3540_));
 sky130_fd_sc_hd__buf_1 _7195_ (.A(_3540_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_2 _7196_ (.A0(\rf.registers[7][21] ),
    .A1(_3500_),
    .S(_3539_),
    .X(_3541_));
 sky130_fd_sc_hd__buf_1 _7197_ (.A(_3541_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_2 _7198_ (.A0(\rf.registers[7][22] ),
    .A1(_3502_),
    .S(_3539_),
    .X(_3542_));
 sky130_fd_sc_hd__buf_1 _7199_ (.A(_3542_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_2 _7200_ (.A0(\rf.registers[7][23] ),
    .A1(_3504_),
    .S(_3539_),
    .X(_3543_));
 sky130_fd_sc_hd__buf_1 _7201_ (.A(_3543_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_2 _7202_ (.A0(\rf.registers[7][24] ),
    .A1(_3506_),
    .S(_3539_),
    .X(_3544_));
 sky130_fd_sc_hd__buf_1 _7203_ (.A(_3544_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_2 _7204_ (.A0(\rf.registers[7][25] ),
    .A1(_3508_),
    .S(_3539_),
    .X(_3545_));
 sky130_fd_sc_hd__buf_1 _7205_ (.A(_3545_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_2 _7206_ (.A0(\rf.registers[7][26] ),
    .A1(_3442_),
    .S(_3539_),
    .X(_3546_));
 sky130_fd_sc_hd__buf_1 _7207_ (.A(_3546_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_2 _7208_ (.A0(\rf.registers[7][27] ),
    .A1(_3444_),
    .S(_3539_),
    .X(_3547_));
 sky130_fd_sc_hd__buf_1 _7209_ (.A(_3547_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_2 _7210_ (.A0(\rf.registers[7][28] ),
    .A1(_3446_),
    .S(_3539_),
    .X(_3548_));
 sky130_fd_sc_hd__buf_1 _7211_ (.A(_3548_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_2 _7212_ (.A0(\rf.registers[7][29] ),
    .A1(_3448_),
    .S(_3539_),
    .X(_3549_));
 sky130_fd_sc_hd__buf_1 _7213_ (.A(_3549_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_2 _7214_ (.A0(\rf.registers[7][30] ),
    .A1(_3450_),
    .S(_3516_),
    .X(_3550_));
 sky130_fd_sc_hd__buf_1 _7215_ (.A(_3550_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_2 _7216_ (.A0(\rf.registers[7][31] ),
    .A1(_3452_),
    .S(_3516_),
    .X(_3551_));
 sky130_fd_sc_hd__buf_1 _7217_ (.A(_3551_),
    .X(_0117_));
 sky130_fd_sc_hd__and3b_2 _7218_ (.A_N(A3[1]),
    .B(A3[0]),
    .C(WE3),
    .X(_3552_));
 sky130_fd_sc_hd__and3_2 _7219_ (.A(A3[4]),
    .B(A3[3]),
    .C(A3[2]),
    .X(_3553_));
 sky130_fd_sc_hd__nand2_2 _7220_ (.A(_3552_),
    .B(_3553_),
    .Y(_3554_));
 sky130_fd_sc_hd__buf_1 _7221_ (.A(_3554_),
    .X(_3555_));
 sky130_fd_sc_hd__mux2_2 _7222_ (.A0(_3019_),
    .A1(\rf.registers[29][0] ),
    .S(_3555_),
    .X(_3556_));
 sky130_fd_sc_hd__buf_1 _7223_ (.A(_3556_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_2 _7224_ (.A0(_3025_),
    .A1(\rf.registers[29][1] ),
    .S(_3555_),
    .X(_3557_));
 sky130_fd_sc_hd__buf_1 _7225_ (.A(_3557_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_2 _7226_ (.A0(_3027_),
    .A1(\rf.registers[29][2] ),
    .S(_3555_),
    .X(_3558_));
 sky130_fd_sc_hd__buf_1 _7227_ (.A(_3558_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_2 _7228_ (.A0(_3029_),
    .A1(\rf.registers[29][3] ),
    .S(_3555_),
    .X(_3559_));
 sky130_fd_sc_hd__buf_1 _7229_ (.A(_3559_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_2 _7230_ (.A0(_3031_),
    .A1(\rf.registers[29][4] ),
    .S(_3555_),
    .X(_3560_));
 sky130_fd_sc_hd__buf_1 _7231_ (.A(_3560_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_2 _7232_ (.A0(_3033_),
    .A1(\rf.registers[29][5] ),
    .S(_3555_),
    .X(_3561_));
 sky130_fd_sc_hd__buf_1 _7233_ (.A(_3561_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_2 _7234_ (.A0(_3035_),
    .A1(\rf.registers[29][6] ),
    .S(_3555_),
    .X(_3562_));
 sky130_fd_sc_hd__buf_1 _7235_ (.A(_3562_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_2 _7236_ (.A0(_3037_),
    .A1(\rf.registers[29][7] ),
    .S(_3555_),
    .X(_3563_));
 sky130_fd_sc_hd__buf_1 _7237_ (.A(_3563_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_2 _7238_ (.A0(_3039_),
    .A1(\rf.registers[29][8] ),
    .S(_3555_),
    .X(_3564_));
 sky130_fd_sc_hd__buf_1 _7239_ (.A(_3564_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_2 _7240_ (.A0(_3041_),
    .A1(\rf.registers[29][9] ),
    .S(_3555_),
    .X(_3565_));
 sky130_fd_sc_hd__buf_1 _7241_ (.A(_3565_),
    .X(_0127_));
 sky130_fd_sc_hd__buf_1 _7242_ (.A(_3554_),
    .X(_3566_));
 sky130_fd_sc_hd__mux2_2 _7243_ (.A0(_3043_),
    .A1(\rf.registers[29][10] ),
    .S(_3566_),
    .X(_3567_));
 sky130_fd_sc_hd__buf_1 _7244_ (.A(_3567_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_2 _7245_ (.A0(_3046_),
    .A1(\rf.registers[29][11] ),
    .S(_3566_),
    .X(_3568_));
 sky130_fd_sc_hd__buf_1 _7246_ (.A(_3568_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_2 _7247_ (.A0(_3048_),
    .A1(\rf.registers[29][12] ),
    .S(_3566_),
    .X(_3569_));
 sky130_fd_sc_hd__buf_1 _7248_ (.A(_3569_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_2 _7249_ (.A0(_3050_),
    .A1(\rf.registers[29][13] ),
    .S(_3566_),
    .X(_3570_));
 sky130_fd_sc_hd__buf_1 _7250_ (.A(_3570_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_2 _7251_ (.A0(_3052_),
    .A1(\rf.registers[29][14] ),
    .S(_3566_),
    .X(_3571_));
 sky130_fd_sc_hd__buf_1 _7252_ (.A(_3571_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_2 _7253_ (.A0(_3054_),
    .A1(\rf.registers[29][15] ),
    .S(_3566_),
    .X(_3572_));
 sky130_fd_sc_hd__buf_1 _7254_ (.A(_3572_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_2 _7255_ (.A0(_3056_),
    .A1(\rf.registers[29][16] ),
    .S(_3566_),
    .X(_3573_));
 sky130_fd_sc_hd__buf_1 _7256_ (.A(_3573_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_2 _7257_ (.A0(_3058_),
    .A1(\rf.registers[29][17] ),
    .S(_3566_),
    .X(_3574_));
 sky130_fd_sc_hd__buf_1 _7258_ (.A(_3574_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_2 _7259_ (.A0(_3060_),
    .A1(\rf.registers[29][18] ),
    .S(_3566_),
    .X(_3575_));
 sky130_fd_sc_hd__buf_1 _7260_ (.A(_3575_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_2 _7261_ (.A0(_3062_),
    .A1(\rf.registers[29][19] ),
    .S(_3566_),
    .X(_3576_));
 sky130_fd_sc_hd__buf_1 _7262_ (.A(_3576_),
    .X(_0137_));
 sky130_fd_sc_hd__buf_1 _7263_ (.A(_3554_),
    .X(_3577_));
 sky130_fd_sc_hd__mux2_2 _7264_ (.A0(_3064_),
    .A1(\rf.registers[29][20] ),
    .S(_3577_),
    .X(_3578_));
 sky130_fd_sc_hd__buf_1 _7265_ (.A(_3578_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_2 _7266_ (.A0(_3067_),
    .A1(\rf.registers[29][21] ),
    .S(_3577_),
    .X(_3579_));
 sky130_fd_sc_hd__buf_1 _7267_ (.A(_3579_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_2 _7268_ (.A0(_3069_),
    .A1(\rf.registers[29][22] ),
    .S(_3577_),
    .X(_3580_));
 sky130_fd_sc_hd__buf_1 _7269_ (.A(_3580_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_2 _7270_ (.A0(_3071_),
    .A1(\rf.registers[29][23] ),
    .S(_3577_),
    .X(_3581_));
 sky130_fd_sc_hd__buf_1 _7271_ (.A(_3581_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_2 _7272_ (.A0(_3073_),
    .A1(\rf.registers[29][24] ),
    .S(_3577_),
    .X(_3582_));
 sky130_fd_sc_hd__buf_1 _7273_ (.A(_3582_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_2 _7274_ (.A0(_3075_),
    .A1(\rf.registers[29][25] ),
    .S(_3577_),
    .X(_3583_));
 sky130_fd_sc_hd__buf_1 _7275_ (.A(_3583_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_2 _7276_ (.A0(_3077_),
    .A1(\rf.registers[29][26] ),
    .S(_3577_),
    .X(_3584_));
 sky130_fd_sc_hd__buf_1 _7277_ (.A(_3584_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_2 _7278_ (.A0(_3079_),
    .A1(\rf.registers[29][27] ),
    .S(_3577_),
    .X(_3585_));
 sky130_fd_sc_hd__buf_1 _7279_ (.A(_3585_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_2 _7280_ (.A0(_3081_),
    .A1(\rf.registers[29][28] ),
    .S(_3577_),
    .X(_3586_));
 sky130_fd_sc_hd__buf_1 _7281_ (.A(_3586_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_2 _7282_ (.A0(_3083_),
    .A1(\rf.registers[29][29] ),
    .S(_3577_),
    .X(_3587_));
 sky130_fd_sc_hd__buf_1 _7283_ (.A(_3587_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_2 _7284_ (.A0(_3085_),
    .A1(\rf.registers[29][30] ),
    .S(_3554_),
    .X(_3588_));
 sky130_fd_sc_hd__buf_1 _7285_ (.A(_3588_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_2 _7286_ (.A0(_3087_),
    .A1(\rf.registers[29][31] ),
    .S(_3554_),
    .X(_3589_));
 sky130_fd_sc_hd__buf_1 _7287_ (.A(_3589_),
    .X(_0149_));
 sky130_fd_sc_hd__nand2_2 _7288_ (.A(_3193_),
    .B(_3553_),
    .Y(_3590_));
 sky130_fd_sc_hd__buf_1 _7289_ (.A(_3590_),
    .X(_3591_));
 sky130_fd_sc_hd__mux2_2 _7290_ (.A0(_3019_),
    .A1(\rf.registers[31][0] ),
    .S(_3591_),
    .X(_3592_));
 sky130_fd_sc_hd__buf_1 _7291_ (.A(_3592_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_2 _7292_ (.A0(_3025_),
    .A1(\rf.registers[31][1] ),
    .S(_3591_),
    .X(_3593_));
 sky130_fd_sc_hd__buf_1 _7293_ (.A(_3593_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_2 _7294_ (.A0(_3027_),
    .A1(\rf.registers[31][2] ),
    .S(_3591_),
    .X(_3594_));
 sky130_fd_sc_hd__buf_1 _7295_ (.A(_3594_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_2 _7296_ (.A0(_3029_),
    .A1(\rf.registers[31][3] ),
    .S(_3591_),
    .X(_3595_));
 sky130_fd_sc_hd__buf_1 _7297_ (.A(_3595_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_2 _7298_ (.A0(_3031_),
    .A1(\rf.registers[31][4] ),
    .S(_3591_),
    .X(_3596_));
 sky130_fd_sc_hd__buf_1 _7299_ (.A(_3596_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_2 _7300_ (.A0(_3033_),
    .A1(\rf.registers[31][5] ),
    .S(_3591_),
    .X(_3597_));
 sky130_fd_sc_hd__buf_1 _7301_ (.A(_3597_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_2 _7302_ (.A0(_3035_),
    .A1(\rf.registers[31][6] ),
    .S(_3591_),
    .X(_3598_));
 sky130_fd_sc_hd__buf_1 _7303_ (.A(_3598_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_2 _7304_ (.A0(_3037_),
    .A1(\rf.registers[31][7] ),
    .S(_3591_),
    .X(_3599_));
 sky130_fd_sc_hd__buf_1 _7305_ (.A(_3599_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_2 _7306_ (.A0(_3039_),
    .A1(\rf.registers[31][8] ),
    .S(_3591_),
    .X(_3600_));
 sky130_fd_sc_hd__buf_1 _7307_ (.A(_3600_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_2 _7308_ (.A0(_3041_),
    .A1(\rf.registers[31][9] ),
    .S(_3591_),
    .X(_3601_));
 sky130_fd_sc_hd__buf_1 _7309_ (.A(_3601_),
    .X(_0159_));
 sky130_fd_sc_hd__buf_1 _7310_ (.A(_3590_),
    .X(_3602_));
 sky130_fd_sc_hd__mux2_2 _7311_ (.A0(_3043_),
    .A1(\rf.registers[31][10] ),
    .S(_3602_),
    .X(_3603_));
 sky130_fd_sc_hd__buf_1 _7312_ (.A(_3603_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_2 _7313_ (.A0(_3046_),
    .A1(\rf.registers[31][11] ),
    .S(_3602_),
    .X(_3604_));
 sky130_fd_sc_hd__buf_1 _7314_ (.A(_3604_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_2 _7315_ (.A0(_3048_),
    .A1(\rf.registers[31][12] ),
    .S(_3602_),
    .X(_3605_));
 sky130_fd_sc_hd__buf_1 _7316_ (.A(_3605_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_2 _7317_ (.A0(_3050_),
    .A1(\rf.registers[31][13] ),
    .S(_3602_),
    .X(_3606_));
 sky130_fd_sc_hd__buf_1 _7318_ (.A(_3606_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_2 _7319_ (.A0(_3052_),
    .A1(\rf.registers[31][14] ),
    .S(_3602_),
    .X(_3607_));
 sky130_fd_sc_hd__buf_1 _7320_ (.A(_3607_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_2 _7321_ (.A0(_3054_),
    .A1(\rf.registers[31][15] ),
    .S(_3602_),
    .X(_3608_));
 sky130_fd_sc_hd__buf_1 _7322_ (.A(_3608_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_2 _7323_ (.A0(_3056_),
    .A1(\rf.registers[31][16] ),
    .S(_3602_),
    .X(_3609_));
 sky130_fd_sc_hd__buf_1 _7324_ (.A(_3609_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_2 _7325_ (.A0(_3058_),
    .A1(\rf.registers[31][17] ),
    .S(_3602_),
    .X(_3610_));
 sky130_fd_sc_hd__buf_1 _7326_ (.A(_3610_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_2 _7327_ (.A0(_3060_),
    .A1(\rf.registers[31][18] ),
    .S(_3602_),
    .X(_3611_));
 sky130_fd_sc_hd__buf_1 _7328_ (.A(_3611_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_2 _7329_ (.A0(_3062_),
    .A1(\rf.registers[31][19] ),
    .S(_3602_),
    .X(_3612_));
 sky130_fd_sc_hd__buf_1 _7330_ (.A(_3612_),
    .X(_0169_));
 sky130_fd_sc_hd__buf_1 _7331_ (.A(_3590_),
    .X(_3613_));
 sky130_fd_sc_hd__mux2_2 _7332_ (.A0(_3064_),
    .A1(\rf.registers[31][20] ),
    .S(_3613_),
    .X(_3614_));
 sky130_fd_sc_hd__buf_1 _7333_ (.A(_3614_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_2 _7334_ (.A0(_3067_),
    .A1(\rf.registers[31][21] ),
    .S(_3613_),
    .X(_3615_));
 sky130_fd_sc_hd__buf_1 _7335_ (.A(_3615_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_2 _7336_ (.A0(_3069_),
    .A1(\rf.registers[31][22] ),
    .S(_3613_),
    .X(_3616_));
 sky130_fd_sc_hd__buf_1 _7337_ (.A(_3616_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_2 _7338_ (.A0(_3071_),
    .A1(\rf.registers[31][23] ),
    .S(_3613_),
    .X(_3617_));
 sky130_fd_sc_hd__buf_1 _7339_ (.A(_3617_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_2 _7340_ (.A0(_3073_),
    .A1(\rf.registers[31][24] ),
    .S(_3613_),
    .X(_3618_));
 sky130_fd_sc_hd__buf_1 _7341_ (.A(_3618_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_2 _7342_ (.A0(_3075_),
    .A1(\rf.registers[31][25] ),
    .S(_3613_),
    .X(_3619_));
 sky130_fd_sc_hd__buf_1 _7343_ (.A(_3619_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_2 _7344_ (.A0(_3077_),
    .A1(\rf.registers[31][26] ),
    .S(_3613_),
    .X(_3620_));
 sky130_fd_sc_hd__buf_1 _7345_ (.A(_3620_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_2 _7346_ (.A0(_3079_),
    .A1(\rf.registers[31][27] ),
    .S(_3613_),
    .X(_3621_));
 sky130_fd_sc_hd__buf_1 _7347_ (.A(_3621_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_2 _7348_ (.A0(_3081_),
    .A1(\rf.registers[31][28] ),
    .S(_3613_),
    .X(_3622_));
 sky130_fd_sc_hd__buf_1 _7349_ (.A(_3622_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_2 _7350_ (.A0(_3083_),
    .A1(\rf.registers[31][29] ),
    .S(_3613_),
    .X(_3623_));
 sky130_fd_sc_hd__buf_1 _7351_ (.A(_3623_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_2 _7352_ (.A0(_3085_),
    .A1(\rf.registers[31][30] ),
    .S(_3590_),
    .X(_3624_));
 sky130_fd_sc_hd__buf_1 _7353_ (.A(_3624_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_2 _7354_ (.A0(_3087_),
    .A1(\rf.registers[31][31] ),
    .S(_3590_),
    .X(_3625_));
 sky130_fd_sc_hd__buf_1 _7355_ (.A(_3625_),
    .X(_0181_));
 sky130_fd_sc_hd__and3b_2 _7356_ (.A_N(A3[2]),
    .B(A3[3]),
    .C(A3[4]),
    .X(_3626_));
 sky130_fd_sc_hd__nand2_2 _7357_ (.A(_3020_),
    .B(_3626_),
    .Y(_3627_));
 sky130_fd_sc_hd__buf_1 _7358_ (.A(_3627_),
    .X(_3628_));
 sky130_fd_sc_hd__mux2_2 _7359_ (.A0(_3019_),
    .A1(\rf.registers[26][0] ),
    .S(_3628_),
    .X(_3629_));
 sky130_fd_sc_hd__buf_1 _7360_ (.A(_3629_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_2 _7361_ (.A0(_3025_),
    .A1(\rf.registers[26][1] ),
    .S(_3628_),
    .X(_3630_));
 sky130_fd_sc_hd__buf_1 _7362_ (.A(_3630_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_2 _7363_ (.A0(_3027_),
    .A1(\rf.registers[26][2] ),
    .S(_3628_),
    .X(_3631_));
 sky130_fd_sc_hd__buf_1 _7364_ (.A(_3631_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_2 _7365_ (.A0(_3029_),
    .A1(\rf.registers[26][3] ),
    .S(_3628_),
    .X(_3632_));
 sky130_fd_sc_hd__buf_1 _7366_ (.A(_3632_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_2 _7367_ (.A0(_3031_),
    .A1(\rf.registers[26][4] ),
    .S(_3628_),
    .X(_3633_));
 sky130_fd_sc_hd__buf_1 _7368_ (.A(_3633_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_2 _7369_ (.A0(_3033_),
    .A1(\rf.registers[26][5] ),
    .S(_3628_),
    .X(_3634_));
 sky130_fd_sc_hd__buf_1 _7370_ (.A(_3634_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_2 _7371_ (.A0(_3035_),
    .A1(\rf.registers[26][6] ),
    .S(_3628_),
    .X(_3635_));
 sky130_fd_sc_hd__buf_1 _7372_ (.A(_3635_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_2 _7373_ (.A0(_3037_),
    .A1(\rf.registers[26][7] ),
    .S(_3628_),
    .X(_3636_));
 sky130_fd_sc_hd__buf_1 _7374_ (.A(_3636_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_2 _7375_ (.A0(_3039_),
    .A1(\rf.registers[26][8] ),
    .S(_3628_),
    .X(_3637_));
 sky130_fd_sc_hd__buf_1 _7376_ (.A(_3637_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_2 _7377_ (.A0(_3041_),
    .A1(\rf.registers[26][9] ),
    .S(_3628_),
    .X(_3638_));
 sky130_fd_sc_hd__buf_1 _7378_ (.A(_3638_),
    .X(_0191_));
 sky130_fd_sc_hd__buf_1 _7379_ (.A(_3627_),
    .X(_3639_));
 sky130_fd_sc_hd__mux2_2 _7380_ (.A0(_3043_),
    .A1(\rf.registers[26][10] ),
    .S(_3639_),
    .X(_3640_));
 sky130_fd_sc_hd__buf_1 _7381_ (.A(_3640_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_2 _7382_ (.A0(_3046_),
    .A1(\rf.registers[26][11] ),
    .S(_3639_),
    .X(_3641_));
 sky130_fd_sc_hd__buf_1 _7383_ (.A(_3641_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_2 _7384_ (.A0(_3048_),
    .A1(\rf.registers[26][12] ),
    .S(_3639_),
    .X(_3642_));
 sky130_fd_sc_hd__buf_1 _7385_ (.A(_3642_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_2 _7386_ (.A0(_3050_),
    .A1(\rf.registers[26][13] ),
    .S(_3639_),
    .X(_3643_));
 sky130_fd_sc_hd__buf_1 _7387_ (.A(_3643_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_2 _7388_ (.A0(_3052_),
    .A1(\rf.registers[26][14] ),
    .S(_3639_),
    .X(_3644_));
 sky130_fd_sc_hd__buf_1 _7389_ (.A(_3644_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_2 _7390_ (.A0(_3054_),
    .A1(\rf.registers[26][15] ),
    .S(_3639_),
    .X(_3645_));
 sky130_fd_sc_hd__buf_1 _7391_ (.A(_3645_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_2 _7392_ (.A0(_3056_),
    .A1(\rf.registers[26][16] ),
    .S(_3639_),
    .X(_3646_));
 sky130_fd_sc_hd__buf_1 _7393_ (.A(_3646_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_2 _7394_ (.A0(_3058_),
    .A1(\rf.registers[26][17] ),
    .S(_3639_),
    .X(_3647_));
 sky130_fd_sc_hd__buf_1 _7395_ (.A(_3647_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_2 _7396_ (.A0(_3060_),
    .A1(\rf.registers[26][18] ),
    .S(_3639_),
    .X(_3648_));
 sky130_fd_sc_hd__buf_1 _7397_ (.A(_3648_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_2 _7398_ (.A0(_3062_),
    .A1(\rf.registers[26][19] ),
    .S(_3639_),
    .X(_3649_));
 sky130_fd_sc_hd__buf_1 _7399_ (.A(_3649_),
    .X(_0201_));
 sky130_fd_sc_hd__buf_1 _7400_ (.A(_3627_),
    .X(_3650_));
 sky130_fd_sc_hd__mux2_2 _7401_ (.A0(_3064_),
    .A1(\rf.registers[26][20] ),
    .S(_3650_),
    .X(_3651_));
 sky130_fd_sc_hd__buf_1 _7402_ (.A(_3651_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_2 _7403_ (.A0(_3067_),
    .A1(\rf.registers[26][21] ),
    .S(_3650_),
    .X(_3652_));
 sky130_fd_sc_hd__buf_1 _7404_ (.A(_3652_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_2 _7405_ (.A0(_3069_),
    .A1(\rf.registers[26][22] ),
    .S(_3650_),
    .X(_3653_));
 sky130_fd_sc_hd__buf_1 _7406_ (.A(_3653_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_2 _7407_ (.A0(_3071_),
    .A1(\rf.registers[26][23] ),
    .S(_3650_),
    .X(_3654_));
 sky130_fd_sc_hd__buf_1 _7408_ (.A(_3654_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_2 _7409_ (.A0(_3073_),
    .A1(\rf.registers[26][24] ),
    .S(_3650_),
    .X(_3655_));
 sky130_fd_sc_hd__buf_1 _7410_ (.A(_3655_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_2 _7411_ (.A0(_3075_),
    .A1(\rf.registers[26][25] ),
    .S(_3650_),
    .X(_3656_));
 sky130_fd_sc_hd__buf_1 _7412_ (.A(_3656_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_2 _7413_ (.A0(_3077_),
    .A1(\rf.registers[26][26] ),
    .S(_3650_),
    .X(_3657_));
 sky130_fd_sc_hd__buf_1 _7414_ (.A(_3657_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_2 _7415_ (.A0(_3079_),
    .A1(\rf.registers[26][27] ),
    .S(_3650_),
    .X(_3658_));
 sky130_fd_sc_hd__buf_1 _7416_ (.A(_3658_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_2 _7417_ (.A0(_3081_),
    .A1(\rf.registers[26][28] ),
    .S(_3650_),
    .X(_3659_));
 sky130_fd_sc_hd__buf_1 _7418_ (.A(_3659_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_2 _7419_ (.A0(_3083_),
    .A1(\rf.registers[26][29] ),
    .S(_3650_),
    .X(_3660_));
 sky130_fd_sc_hd__buf_1 _7420_ (.A(_3660_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_2 _7421_ (.A0(_3085_),
    .A1(\rf.registers[26][30] ),
    .S(_3627_),
    .X(_3661_));
 sky130_fd_sc_hd__buf_1 _7422_ (.A(_3661_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_2 _7423_ (.A0(_3087_),
    .A1(\rf.registers[26][31] ),
    .S(_3627_),
    .X(_3662_));
 sky130_fd_sc_hd__buf_1 _7424_ (.A(_3662_),
    .X(_0213_));
 sky130_fd_sc_hd__nand2_2 _7425_ (.A(_3552_),
    .B(_3626_),
    .Y(_3663_));
 sky130_fd_sc_hd__buf_1 _7426_ (.A(_3663_),
    .X(_3664_));
 sky130_fd_sc_hd__mux2_2 _7427_ (.A0(_3019_),
    .A1(\rf.registers[25][0] ),
    .S(_3664_),
    .X(_3665_));
 sky130_fd_sc_hd__buf_1 _7428_ (.A(_3665_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_2 _7429_ (.A0(_3025_),
    .A1(\rf.registers[25][1] ),
    .S(_3664_),
    .X(_3666_));
 sky130_fd_sc_hd__buf_1 _7430_ (.A(_3666_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_2 _7431_ (.A0(_3027_),
    .A1(\rf.registers[25][2] ),
    .S(_3664_),
    .X(_3667_));
 sky130_fd_sc_hd__buf_1 _7432_ (.A(_3667_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_2 _7433_ (.A0(_3029_),
    .A1(\rf.registers[25][3] ),
    .S(_3664_),
    .X(_3668_));
 sky130_fd_sc_hd__buf_1 _7434_ (.A(_3668_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_2 _7435_ (.A0(_3031_),
    .A1(\rf.registers[25][4] ),
    .S(_3664_),
    .X(_3669_));
 sky130_fd_sc_hd__buf_1 _7436_ (.A(_3669_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_2 _7437_ (.A0(_3033_),
    .A1(\rf.registers[25][5] ),
    .S(_3664_),
    .X(_3670_));
 sky130_fd_sc_hd__buf_1 _7438_ (.A(_3670_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_2 _7439_ (.A0(_3035_),
    .A1(\rf.registers[25][6] ),
    .S(_3664_),
    .X(_3671_));
 sky130_fd_sc_hd__buf_1 _7440_ (.A(_3671_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_2 _7441_ (.A0(_3037_),
    .A1(\rf.registers[25][7] ),
    .S(_3664_),
    .X(_3672_));
 sky130_fd_sc_hd__buf_1 _7442_ (.A(_3672_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_2 _7443_ (.A0(_3039_),
    .A1(\rf.registers[25][8] ),
    .S(_3664_),
    .X(_3673_));
 sky130_fd_sc_hd__buf_1 _7444_ (.A(_3673_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_2 _7445_ (.A0(_3041_),
    .A1(\rf.registers[25][9] ),
    .S(_3664_),
    .X(_3674_));
 sky130_fd_sc_hd__buf_1 _7446_ (.A(_3674_),
    .X(_0223_));
 sky130_fd_sc_hd__buf_1 _7447_ (.A(_3663_),
    .X(_3675_));
 sky130_fd_sc_hd__mux2_2 _7448_ (.A0(_3043_),
    .A1(\rf.registers[25][10] ),
    .S(_3675_),
    .X(_3676_));
 sky130_fd_sc_hd__buf_1 _7449_ (.A(_3676_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_2 _7450_ (.A0(_3046_),
    .A1(\rf.registers[25][11] ),
    .S(_3675_),
    .X(_3677_));
 sky130_fd_sc_hd__buf_1 _7451_ (.A(_3677_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_2 _7452_ (.A0(_3048_),
    .A1(\rf.registers[25][12] ),
    .S(_3675_),
    .X(_3678_));
 sky130_fd_sc_hd__buf_1 _7453_ (.A(_3678_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_2 _7454_ (.A0(_3050_),
    .A1(\rf.registers[25][13] ),
    .S(_3675_),
    .X(_3679_));
 sky130_fd_sc_hd__buf_1 _7455_ (.A(_3679_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_2 _7456_ (.A0(_3052_),
    .A1(\rf.registers[25][14] ),
    .S(_3675_),
    .X(_3680_));
 sky130_fd_sc_hd__buf_1 _7457_ (.A(_3680_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_2 _7458_ (.A0(_3054_),
    .A1(\rf.registers[25][15] ),
    .S(_3675_),
    .X(_3681_));
 sky130_fd_sc_hd__buf_1 _7459_ (.A(_3681_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_2 _7460_ (.A0(_3056_),
    .A1(\rf.registers[25][16] ),
    .S(_3675_),
    .X(_3682_));
 sky130_fd_sc_hd__buf_1 _7461_ (.A(_3682_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_2 _7462_ (.A0(_3058_),
    .A1(\rf.registers[25][17] ),
    .S(_3675_),
    .X(_3683_));
 sky130_fd_sc_hd__buf_1 _7463_ (.A(_3683_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_2 _7464_ (.A0(_3060_),
    .A1(\rf.registers[25][18] ),
    .S(_3675_),
    .X(_3684_));
 sky130_fd_sc_hd__buf_1 _7465_ (.A(_3684_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_2 _7466_ (.A0(_3062_),
    .A1(\rf.registers[25][19] ),
    .S(_3675_),
    .X(_3685_));
 sky130_fd_sc_hd__buf_1 _7467_ (.A(_3685_),
    .X(_0233_));
 sky130_fd_sc_hd__buf_1 _7468_ (.A(_3663_),
    .X(_3686_));
 sky130_fd_sc_hd__mux2_2 _7469_ (.A0(_3064_),
    .A1(\rf.registers[25][20] ),
    .S(_3686_),
    .X(_3687_));
 sky130_fd_sc_hd__buf_1 _7470_ (.A(_3687_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_2 _7471_ (.A0(_3067_),
    .A1(\rf.registers[25][21] ),
    .S(_3686_),
    .X(_3688_));
 sky130_fd_sc_hd__buf_1 _7472_ (.A(_3688_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_2 _7473_ (.A0(_3069_),
    .A1(\rf.registers[25][22] ),
    .S(_3686_),
    .X(_3689_));
 sky130_fd_sc_hd__buf_1 _7474_ (.A(_3689_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_2 _7475_ (.A0(_3071_),
    .A1(\rf.registers[25][23] ),
    .S(_3686_),
    .X(_3690_));
 sky130_fd_sc_hd__buf_1 _7476_ (.A(_3690_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_2 _7477_ (.A0(_3073_),
    .A1(\rf.registers[25][24] ),
    .S(_3686_),
    .X(_3691_));
 sky130_fd_sc_hd__buf_1 _7478_ (.A(_3691_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_2 _7479_ (.A0(_3075_),
    .A1(\rf.registers[25][25] ),
    .S(_3686_),
    .X(_3692_));
 sky130_fd_sc_hd__buf_1 _7480_ (.A(_3692_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_2 _7481_ (.A0(_3077_),
    .A1(\rf.registers[25][26] ),
    .S(_3686_),
    .X(_3693_));
 sky130_fd_sc_hd__buf_1 _7482_ (.A(_3693_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_2 _7483_ (.A0(_3079_),
    .A1(\rf.registers[25][27] ),
    .S(_3686_),
    .X(_3694_));
 sky130_fd_sc_hd__buf_1 _7484_ (.A(_3694_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_2 _7485_ (.A0(_3081_),
    .A1(\rf.registers[25][28] ),
    .S(_3686_),
    .X(_3695_));
 sky130_fd_sc_hd__buf_1 _7486_ (.A(_3695_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_2 _7487_ (.A0(_3083_),
    .A1(\rf.registers[25][29] ),
    .S(_3686_),
    .X(_3696_));
 sky130_fd_sc_hd__buf_1 _7488_ (.A(_3696_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_2 _7489_ (.A0(_3085_),
    .A1(\rf.registers[25][30] ),
    .S(_3663_),
    .X(_3697_));
 sky130_fd_sc_hd__buf_1 _7490_ (.A(_3697_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_2 _7491_ (.A0(_3087_),
    .A1(\rf.registers[25][31] ),
    .S(_3663_),
    .X(_3698_));
 sky130_fd_sc_hd__buf_1 _7492_ (.A(_3698_),
    .X(_0245_));
 sky130_fd_sc_hd__nand2_2 _7493_ (.A(_3193_),
    .B(_3626_),
    .Y(_3699_));
 sky130_fd_sc_hd__buf_1 _7494_ (.A(_3699_),
    .X(_3700_));
 sky130_fd_sc_hd__mux2_2 _7495_ (.A0(_3019_),
    .A1(\rf.registers[27][0] ),
    .S(_3700_),
    .X(_3701_));
 sky130_fd_sc_hd__buf_1 _7496_ (.A(_3701_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_2 _7497_ (.A0(_3025_),
    .A1(\rf.registers[27][1] ),
    .S(_3700_),
    .X(_3702_));
 sky130_fd_sc_hd__buf_1 _7498_ (.A(_3702_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_2 _7499_ (.A0(_3027_),
    .A1(\rf.registers[27][2] ),
    .S(_3700_),
    .X(_3703_));
 sky130_fd_sc_hd__buf_1 _7500_ (.A(_3703_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_2 _7501_ (.A0(_3029_),
    .A1(\rf.registers[27][3] ),
    .S(_3700_),
    .X(_3704_));
 sky130_fd_sc_hd__buf_1 _7502_ (.A(_3704_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_2 _7503_ (.A0(_3031_),
    .A1(\rf.registers[27][4] ),
    .S(_3700_),
    .X(_3705_));
 sky130_fd_sc_hd__buf_1 _7504_ (.A(_3705_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_2 _7505_ (.A0(_3033_),
    .A1(\rf.registers[27][5] ),
    .S(_3700_),
    .X(_3706_));
 sky130_fd_sc_hd__buf_1 _7506_ (.A(_3706_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_2 _7507_ (.A0(_3035_),
    .A1(\rf.registers[27][6] ),
    .S(_3700_),
    .X(_3707_));
 sky130_fd_sc_hd__buf_1 _7508_ (.A(_3707_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_2 _7509_ (.A0(_3037_),
    .A1(\rf.registers[27][7] ),
    .S(_3700_),
    .X(_3708_));
 sky130_fd_sc_hd__buf_1 _7510_ (.A(_3708_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_2 _7511_ (.A0(_3039_),
    .A1(\rf.registers[27][8] ),
    .S(_3700_),
    .X(_3709_));
 sky130_fd_sc_hd__buf_1 _7512_ (.A(_3709_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_2 _7513_ (.A0(_3041_),
    .A1(\rf.registers[27][9] ),
    .S(_3700_),
    .X(_3710_));
 sky130_fd_sc_hd__buf_1 _7514_ (.A(_3710_),
    .X(_0255_));
 sky130_fd_sc_hd__buf_1 _7515_ (.A(_3699_),
    .X(_3711_));
 sky130_fd_sc_hd__mux2_2 _7516_ (.A0(_3043_),
    .A1(\rf.registers[27][10] ),
    .S(_3711_),
    .X(_3712_));
 sky130_fd_sc_hd__buf_1 _7517_ (.A(_3712_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_2 _7518_ (.A0(_3046_),
    .A1(\rf.registers[27][11] ),
    .S(_3711_),
    .X(_3713_));
 sky130_fd_sc_hd__buf_1 _7519_ (.A(_3713_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_2 _7520_ (.A0(_3048_),
    .A1(\rf.registers[27][12] ),
    .S(_3711_),
    .X(_3714_));
 sky130_fd_sc_hd__buf_1 _7521_ (.A(_3714_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_2 _7522_ (.A0(_3050_),
    .A1(\rf.registers[27][13] ),
    .S(_3711_),
    .X(_3715_));
 sky130_fd_sc_hd__buf_1 _7523_ (.A(_3715_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_2 _7524_ (.A0(_3052_),
    .A1(\rf.registers[27][14] ),
    .S(_3711_),
    .X(_3716_));
 sky130_fd_sc_hd__buf_1 _7525_ (.A(_3716_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_2 _7526_ (.A0(_3054_),
    .A1(\rf.registers[27][15] ),
    .S(_3711_),
    .X(_3717_));
 sky130_fd_sc_hd__buf_1 _7527_ (.A(_3717_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_2 _7528_ (.A0(_3056_),
    .A1(\rf.registers[27][16] ),
    .S(_3711_),
    .X(_3718_));
 sky130_fd_sc_hd__buf_1 _7529_ (.A(_3718_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_2 _7530_ (.A0(_3058_),
    .A1(\rf.registers[27][17] ),
    .S(_3711_),
    .X(_3719_));
 sky130_fd_sc_hd__buf_1 _7531_ (.A(_3719_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_2 _7532_ (.A0(_3060_),
    .A1(\rf.registers[27][18] ),
    .S(_3711_),
    .X(_3720_));
 sky130_fd_sc_hd__buf_1 _7533_ (.A(_3720_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_2 _7534_ (.A0(_3062_),
    .A1(\rf.registers[27][19] ),
    .S(_3711_),
    .X(_3721_));
 sky130_fd_sc_hd__buf_1 _7535_ (.A(_3721_),
    .X(_0265_));
 sky130_fd_sc_hd__buf_1 _7536_ (.A(_3699_),
    .X(_3722_));
 sky130_fd_sc_hd__mux2_2 _7537_ (.A0(_3064_),
    .A1(\rf.registers[27][20] ),
    .S(_3722_),
    .X(_3723_));
 sky130_fd_sc_hd__buf_1 _7538_ (.A(_3723_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_2 _7539_ (.A0(_3067_),
    .A1(\rf.registers[27][21] ),
    .S(_3722_),
    .X(_3724_));
 sky130_fd_sc_hd__buf_1 _7540_ (.A(_3724_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_2 _7541_ (.A0(_3069_),
    .A1(\rf.registers[27][22] ),
    .S(_3722_),
    .X(_3725_));
 sky130_fd_sc_hd__buf_1 _7542_ (.A(_3725_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_2 _7543_ (.A0(_3071_),
    .A1(\rf.registers[27][23] ),
    .S(_3722_),
    .X(_3726_));
 sky130_fd_sc_hd__buf_1 _7544_ (.A(_3726_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_2 _7545_ (.A0(_3073_),
    .A1(\rf.registers[27][24] ),
    .S(_3722_),
    .X(_3727_));
 sky130_fd_sc_hd__buf_1 _7546_ (.A(_3727_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_2 _7547_ (.A0(_3075_),
    .A1(\rf.registers[27][25] ),
    .S(_3722_),
    .X(_3728_));
 sky130_fd_sc_hd__buf_1 _7548_ (.A(_3728_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_2 _7549_ (.A0(_3077_),
    .A1(\rf.registers[27][26] ),
    .S(_3722_),
    .X(_3729_));
 sky130_fd_sc_hd__buf_1 _7550_ (.A(_3729_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_2 _7551_ (.A0(_3079_),
    .A1(\rf.registers[27][27] ),
    .S(_3722_),
    .X(_3730_));
 sky130_fd_sc_hd__buf_1 _7552_ (.A(_3730_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_2 _7553_ (.A0(_3081_),
    .A1(\rf.registers[27][28] ),
    .S(_3722_),
    .X(_3731_));
 sky130_fd_sc_hd__buf_1 _7554_ (.A(_3731_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_2 _7555_ (.A0(_3083_),
    .A1(\rf.registers[27][29] ),
    .S(_3722_),
    .X(_3732_));
 sky130_fd_sc_hd__buf_1 _7556_ (.A(_3732_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_2 _7557_ (.A0(_3085_),
    .A1(\rf.registers[27][30] ),
    .S(_3699_),
    .X(_3733_));
 sky130_fd_sc_hd__buf_1 _7558_ (.A(_3733_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_2 _7559_ (.A0(_3087_),
    .A1(\rf.registers[27][31] ),
    .S(_3699_),
    .X(_3734_));
 sky130_fd_sc_hd__buf_1 _7560_ (.A(_3734_),
    .X(_0277_));
 sky130_fd_sc_hd__nand2b_2 _7561_ (.A_N(_3155_),
    .B(_3553_),
    .Y(_3735_));
 sky130_fd_sc_hd__buf_1 _7562_ (.A(_3735_),
    .X(_3736_));
 sky130_fd_sc_hd__mux2_2 _7563_ (.A0(_3019_),
    .A1(\rf.registers[28][0] ),
    .S(_3736_),
    .X(_3737_));
 sky130_fd_sc_hd__buf_1 _7564_ (.A(_3737_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_2 _7565_ (.A0(_3025_),
    .A1(\rf.registers[28][1] ),
    .S(_3736_),
    .X(_3738_));
 sky130_fd_sc_hd__buf_1 _7566_ (.A(_3738_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_2 _7567_ (.A0(_3027_),
    .A1(\rf.registers[28][2] ),
    .S(_3736_),
    .X(_3739_));
 sky130_fd_sc_hd__buf_1 _7568_ (.A(_3739_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_2 _7569_ (.A0(_3029_),
    .A1(\rf.registers[28][3] ),
    .S(_3736_),
    .X(_3740_));
 sky130_fd_sc_hd__buf_1 _7570_ (.A(_3740_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_2 _7571_ (.A0(_3031_),
    .A1(\rf.registers[28][4] ),
    .S(_3736_),
    .X(_3741_));
 sky130_fd_sc_hd__buf_1 _7572_ (.A(_3741_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_2 _7573_ (.A0(_3033_),
    .A1(\rf.registers[28][5] ),
    .S(_3736_),
    .X(_3742_));
 sky130_fd_sc_hd__buf_1 _7574_ (.A(_3742_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_2 _7575_ (.A0(_3035_),
    .A1(\rf.registers[28][6] ),
    .S(_3736_),
    .X(_3743_));
 sky130_fd_sc_hd__buf_1 _7576_ (.A(_3743_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_2 _7577_ (.A0(_3037_),
    .A1(\rf.registers[28][7] ),
    .S(_3736_),
    .X(_3744_));
 sky130_fd_sc_hd__buf_1 _7578_ (.A(_3744_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_2 _7579_ (.A0(_3039_),
    .A1(\rf.registers[28][8] ),
    .S(_3736_),
    .X(_3745_));
 sky130_fd_sc_hd__buf_1 _7580_ (.A(_3745_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_2 _7581_ (.A0(_3041_),
    .A1(\rf.registers[28][9] ),
    .S(_3736_),
    .X(_3746_));
 sky130_fd_sc_hd__buf_1 _7582_ (.A(_3746_),
    .X(_0287_));
 sky130_fd_sc_hd__buf_1 _7583_ (.A(_3735_),
    .X(_3747_));
 sky130_fd_sc_hd__mux2_2 _7584_ (.A0(_3043_),
    .A1(\rf.registers[28][10] ),
    .S(_3747_),
    .X(_3748_));
 sky130_fd_sc_hd__buf_1 _7585_ (.A(_3748_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_2 _7586_ (.A0(_3046_),
    .A1(\rf.registers[28][11] ),
    .S(_3747_),
    .X(_3749_));
 sky130_fd_sc_hd__buf_1 _7587_ (.A(_3749_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_2 _7588_ (.A0(_3048_),
    .A1(\rf.registers[28][12] ),
    .S(_3747_),
    .X(_3750_));
 sky130_fd_sc_hd__buf_1 _7589_ (.A(_3750_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_2 _7590_ (.A0(_3050_),
    .A1(\rf.registers[28][13] ),
    .S(_3747_),
    .X(_3751_));
 sky130_fd_sc_hd__buf_1 _7591_ (.A(_3751_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_2 _7592_ (.A0(_3052_),
    .A1(\rf.registers[28][14] ),
    .S(_3747_),
    .X(_3752_));
 sky130_fd_sc_hd__buf_1 _7593_ (.A(_3752_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_2 _7594_ (.A0(_3054_),
    .A1(\rf.registers[28][15] ),
    .S(_3747_),
    .X(_3753_));
 sky130_fd_sc_hd__buf_1 _7595_ (.A(_3753_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_2 _7596_ (.A0(_3056_),
    .A1(\rf.registers[28][16] ),
    .S(_3747_),
    .X(_3754_));
 sky130_fd_sc_hd__buf_1 _7597_ (.A(_3754_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_2 _7598_ (.A0(_3058_),
    .A1(\rf.registers[28][17] ),
    .S(_3747_),
    .X(_3755_));
 sky130_fd_sc_hd__buf_1 _7599_ (.A(_3755_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_2 _7600_ (.A0(_3060_),
    .A1(\rf.registers[28][18] ),
    .S(_3747_),
    .X(_3756_));
 sky130_fd_sc_hd__buf_1 _7601_ (.A(_3756_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_2 _7602_ (.A0(_3062_),
    .A1(\rf.registers[28][19] ),
    .S(_3747_),
    .X(_3757_));
 sky130_fd_sc_hd__buf_1 _7603_ (.A(_3757_),
    .X(_0297_));
 sky130_fd_sc_hd__buf_1 _7604_ (.A(_3735_),
    .X(_3758_));
 sky130_fd_sc_hd__mux2_2 _7605_ (.A0(_3064_),
    .A1(\rf.registers[28][20] ),
    .S(_3758_),
    .X(_3759_));
 sky130_fd_sc_hd__buf_1 _7606_ (.A(_3759_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_2 _7607_ (.A0(_3067_),
    .A1(\rf.registers[28][21] ),
    .S(_3758_),
    .X(_3760_));
 sky130_fd_sc_hd__buf_1 _7608_ (.A(_3760_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_2 _7609_ (.A0(_3069_),
    .A1(\rf.registers[28][22] ),
    .S(_3758_),
    .X(_3761_));
 sky130_fd_sc_hd__buf_1 _7610_ (.A(_3761_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_2 _7611_ (.A0(_3071_),
    .A1(\rf.registers[28][23] ),
    .S(_3758_),
    .X(_3762_));
 sky130_fd_sc_hd__buf_1 _7612_ (.A(_3762_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_2 _7613_ (.A0(_3073_),
    .A1(\rf.registers[28][24] ),
    .S(_3758_),
    .X(_3763_));
 sky130_fd_sc_hd__buf_1 _7614_ (.A(_3763_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_2 _7615_ (.A0(_3075_),
    .A1(\rf.registers[28][25] ),
    .S(_3758_),
    .X(_3764_));
 sky130_fd_sc_hd__buf_1 _7616_ (.A(_3764_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_2 _7617_ (.A0(_3077_),
    .A1(\rf.registers[28][26] ),
    .S(_3758_),
    .X(_3765_));
 sky130_fd_sc_hd__buf_1 _7618_ (.A(_3765_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_2 _7619_ (.A0(_3079_),
    .A1(\rf.registers[28][27] ),
    .S(_3758_),
    .X(_3766_));
 sky130_fd_sc_hd__buf_1 _7620_ (.A(_3766_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_2 _7621_ (.A0(_3081_),
    .A1(\rf.registers[28][28] ),
    .S(_3758_),
    .X(_3767_));
 sky130_fd_sc_hd__buf_1 _7622_ (.A(_3767_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_2 _7623_ (.A0(_3083_),
    .A1(\rf.registers[28][29] ),
    .S(_3758_),
    .X(_3768_));
 sky130_fd_sc_hd__buf_1 _7624_ (.A(_3768_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_2 _7625_ (.A0(_3085_),
    .A1(\rf.registers[28][30] ),
    .S(_3735_),
    .X(_3769_));
 sky130_fd_sc_hd__buf_1 _7626_ (.A(_3769_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_2 _7627_ (.A0(_3087_),
    .A1(\rf.registers[28][31] ),
    .S(_3735_),
    .X(_3770_));
 sky130_fd_sc_hd__buf_1 _7628_ (.A(_3770_),
    .X(_0309_));
 sky130_fd_sc_hd__nor2_2 _7629_ (.A(_3005_),
    .B(_3153_),
    .Y(_3771_));
 sky130_fd_sc_hd__buf_1 _7630_ (.A(_3771_),
    .X(_3772_));
 sky130_fd_sc_hd__mux2_2 _7631_ (.A0(\rf.registers[2][0] ),
    .A1(_3454_),
    .S(_3772_),
    .X(_3773_));
 sky130_fd_sc_hd__buf_1 _7632_ (.A(_3773_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_2 _7633_ (.A0(\rf.registers[2][1] ),
    .A1(_3458_),
    .S(_3772_),
    .X(_3774_));
 sky130_fd_sc_hd__buf_1 _7634_ (.A(_3774_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_2 _7635_ (.A0(\rf.registers[2][2] ),
    .A1(_3460_),
    .S(_3772_),
    .X(_3775_));
 sky130_fd_sc_hd__buf_1 _7636_ (.A(_3775_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_2 _7637_ (.A0(\rf.registers[2][3] ),
    .A1(_3462_),
    .S(_3772_),
    .X(_3776_));
 sky130_fd_sc_hd__buf_1 _7638_ (.A(_3776_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_2 _7639_ (.A0(\rf.registers[2][4] ),
    .A1(_3464_),
    .S(_3772_),
    .X(_3777_));
 sky130_fd_sc_hd__buf_1 _7640_ (.A(_3777_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_2 _7641_ (.A0(\rf.registers[2][5] ),
    .A1(_3466_),
    .S(_3772_),
    .X(_3778_));
 sky130_fd_sc_hd__buf_1 _7642_ (.A(_3778_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_2 _7643_ (.A0(\rf.registers[2][6] ),
    .A1(_3468_),
    .S(_3772_),
    .X(_3779_));
 sky130_fd_sc_hd__buf_1 _7644_ (.A(_3779_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_2 _7645_ (.A0(\rf.registers[2][7] ),
    .A1(_3470_),
    .S(_3772_),
    .X(_3780_));
 sky130_fd_sc_hd__buf_1 _7646_ (.A(_3780_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_2 _7647_ (.A0(\rf.registers[2][8] ),
    .A1(_3472_),
    .S(_3772_),
    .X(_3781_));
 sky130_fd_sc_hd__buf_1 _7648_ (.A(_3781_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_2 _7649_ (.A0(\rf.registers[2][9] ),
    .A1(_3474_),
    .S(_3772_),
    .X(_3782_));
 sky130_fd_sc_hd__buf_1 _7650_ (.A(_3782_),
    .X(_0319_));
 sky130_fd_sc_hd__buf_1 _7651_ (.A(_3771_),
    .X(_3783_));
 sky130_fd_sc_hd__mux2_2 _7652_ (.A0(\rf.registers[2][10] ),
    .A1(_3476_),
    .S(_3783_),
    .X(_3784_));
 sky130_fd_sc_hd__buf_1 _7653_ (.A(_3784_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_2 _7654_ (.A0(\rf.registers[2][11] ),
    .A1(_3479_),
    .S(_3783_),
    .X(_3785_));
 sky130_fd_sc_hd__buf_1 _7655_ (.A(_3785_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_2 _7656_ (.A0(\rf.registers[2][12] ),
    .A1(_3481_),
    .S(_3783_),
    .X(_3786_));
 sky130_fd_sc_hd__buf_1 _7657_ (.A(_3786_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_2 _7658_ (.A0(\rf.registers[2][13] ),
    .A1(_3483_),
    .S(_3783_),
    .X(_3787_));
 sky130_fd_sc_hd__buf_1 _7659_ (.A(_3787_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_2 _7660_ (.A0(\rf.registers[2][14] ),
    .A1(_3485_),
    .S(_3783_),
    .X(_3788_));
 sky130_fd_sc_hd__buf_1 _7661_ (.A(_3788_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_2 _7662_ (.A0(\rf.registers[2][15] ),
    .A1(_3487_),
    .S(_3783_),
    .X(_3789_));
 sky130_fd_sc_hd__buf_1 _7663_ (.A(_3789_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_2 _7664_ (.A0(\rf.registers[2][16] ),
    .A1(_3489_),
    .S(_3783_),
    .X(_3790_));
 sky130_fd_sc_hd__buf_1 _7665_ (.A(_3790_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_2 _7666_ (.A0(\rf.registers[2][17] ),
    .A1(_3491_),
    .S(_3783_),
    .X(_3791_));
 sky130_fd_sc_hd__buf_1 _7667_ (.A(_3791_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_2 _7668_ (.A0(\rf.registers[2][18] ),
    .A1(_3493_),
    .S(_3783_),
    .X(_3792_));
 sky130_fd_sc_hd__buf_1 _7669_ (.A(_3792_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_2 _7670_ (.A0(\rf.registers[2][19] ),
    .A1(_3495_),
    .S(_3783_),
    .X(_3793_));
 sky130_fd_sc_hd__buf_1 _7671_ (.A(_3793_),
    .X(_0329_));
 sky130_fd_sc_hd__buf_1 _7672_ (.A(_3771_),
    .X(_3794_));
 sky130_fd_sc_hd__mux2_2 _7673_ (.A0(\rf.registers[2][20] ),
    .A1(_3497_),
    .S(_3794_),
    .X(_3795_));
 sky130_fd_sc_hd__buf_1 _7674_ (.A(_3795_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_2 _7675_ (.A0(\rf.registers[2][21] ),
    .A1(_3500_),
    .S(_3794_),
    .X(_3796_));
 sky130_fd_sc_hd__buf_1 _7676_ (.A(_3796_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_2 _7677_ (.A0(\rf.registers[2][22] ),
    .A1(_3502_),
    .S(_3794_),
    .X(_3797_));
 sky130_fd_sc_hd__buf_1 _7678_ (.A(_3797_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_2 _7679_ (.A0(\rf.registers[2][23] ),
    .A1(_3504_),
    .S(_3794_),
    .X(_3798_));
 sky130_fd_sc_hd__buf_1 _7680_ (.A(_3798_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_2 _7681_ (.A0(\rf.registers[2][24] ),
    .A1(_3506_),
    .S(_3794_),
    .X(_3799_));
 sky130_fd_sc_hd__buf_1 _7682_ (.A(_3799_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_2 _7683_ (.A0(\rf.registers[2][25] ),
    .A1(_3508_),
    .S(_3794_),
    .X(_3800_));
 sky130_fd_sc_hd__buf_1 _7684_ (.A(_3800_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_2 _7685_ (.A0(\rf.registers[2][26] ),
    .A1(_3442_),
    .S(_3794_),
    .X(_3801_));
 sky130_fd_sc_hd__buf_1 _7686_ (.A(_3801_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_2 _7687_ (.A0(\rf.registers[2][27] ),
    .A1(_3444_),
    .S(_3794_),
    .X(_3802_));
 sky130_fd_sc_hd__buf_1 _7688_ (.A(_3802_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_2 _7689_ (.A0(\rf.registers[2][28] ),
    .A1(_3446_),
    .S(_3794_),
    .X(_3803_));
 sky130_fd_sc_hd__buf_1 _7690_ (.A(_3803_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_2 _7691_ (.A0(\rf.registers[2][29] ),
    .A1(_3448_),
    .S(_3794_),
    .X(_3804_));
 sky130_fd_sc_hd__buf_1 _7692_ (.A(_3804_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_2 _7693_ (.A0(\rf.registers[2][30] ),
    .A1(_3450_),
    .S(_3771_),
    .X(_3805_));
 sky130_fd_sc_hd__buf_1 _7694_ (.A(_3805_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_2 _7695_ (.A0(\rf.registers[2][31] ),
    .A1(_3452_),
    .S(_3771_),
    .X(_3806_));
 sky130_fd_sc_hd__buf_1 _7696_ (.A(_3806_),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_2 _7697_ (.A(_3020_),
    .B(_3553_),
    .Y(_3807_));
 sky130_fd_sc_hd__buf_1 _7698_ (.A(_3807_),
    .X(_3808_));
 sky130_fd_sc_hd__mux2_2 _7699_ (.A0(_3019_),
    .A1(\rf.registers[30][0] ),
    .S(_3808_),
    .X(_3809_));
 sky130_fd_sc_hd__buf_1 _7700_ (.A(_3809_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_2 _7701_ (.A0(_3025_),
    .A1(\rf.registers[30][1] ),
    .S(_3808_),
    .X(_3810_));
 sky130_fd_sc_hd__buf_1 _7702_ (.A(_3810_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_2 _7703_ (.A0(_3027_),
    .A1(\rf.registers[30][2] ),
    .S(_3808_),
    .X(_3811_));
 sky130_fd_sc_hd__buf_1 _7704_ (.A(_3811_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_2 _7705_ (.A0(_3029_),
    .A1(\rf.registers[30][3] ),
    .S(_3808_),
    .X(_3812_));
 sky130_fd_sc_hd__buf_1 _7706_ (.A(_3812_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_2 _7707_ (.A0(_3031_),
    .A1(\rf.registers[30][4] ),
    .S(_3808_),
    .X(_3813_));
 sky130_fd_sc_hd__buf_1 _7708_ (.A(_3813_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_2 _7709_ (.A0(_3033_),
    .A1(\rf.registers[30][5] ),
    .S(_3808_),
    .X(_3814_));
 sky130_fd_sc_hd__buf_1 _7710_ (.A(_3814_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_2 _7711_ (.A0(_3035_),
    .A1(\rf.registers[30][6] ),
    .S(_3808_),
    .X(_3815_));
 sky130_fd_sc_hd__buf_1 _7712_ (.A(_3815_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_2 _7713_ (.A0(_3037_),
    .A1(\rf.registers[30][7] ),
    .S(_3808_),
    .X(_3816_));
 sky130_fd_sc_hd__buf_1 _7714_ (.A(_3816_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_2 _7715_ (.A0(_3039_),
    .A1(\rf.registers[30][8] ),
    .S(_3808_),
    .X(_3817_));
 sky130_fd_sc_hd__buf_1 _7716_ (.A(_3817_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_2 _7717_ (.A0(_3041_),
    .A1(\rf.registers[30][9] ),
    .S(_3808_),
    .X(_3818_));
 sky130_fd_sc_hd__buf_1 _7718_ (.A(_3818_),
    .X(_0351_));
 sky130_fd_sc_hd__buf_1 _7719_ (.A(_3807_),
    .X(_3819_));
 sky130_fd_sc_hd__mux2_2 _7720_ (.A0(_3043_),
    .A1(\rf.registers[30][10] ),
    .S(_3819_),
    .X(_3820_));
 sky130_fd_sc_hd__buf_1 _7721_ (.A(_3820_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_2 _7722_ (.A0(_3046_),
    .A1(\rf.registers[30][11] ),
    .S(_3819_),
    .X(_3821_));
 sky130_fd_sc_hd__buf_1 _7723_ (.A(_3821_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_2 _7724_ (.A0(_3048_),
    .A1(\rf.registers[30][12] ),
    .S(_3819_),
    .X(_3822_));
 sky130_fd_sc_hd__buf_1 _7725_ (.A(_3822_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_2 _7726_ (.A0(_3050_),
    .A1(\rf.registers[30][13] ),
    .S(_3819_),
    .X(_3823_));
 sky130_fd_sc_hd__buf_1 _7727_ (.A(_3823_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_2 _7728_ (.A0(_3052_),
    .A1(\rf.registers[30][14] ),
    .S(_3819_),
    .X(_3824_));
 sky130_fd_sc_hd__buf_1 _7729_ (.A(_3824_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_2 _7730_ (.A0(_3054_),
    .A1(\rf.registers[30][15] ),
    .S(_3819_),
    .X(_3825_));
 sky130_fd_sc_hd__buf_1 _7731_ (.A(_3825_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_2 _7732_ (.A0(_3056_),
    .A1(\rf.registers[30][16] ),
    .S(_3819_),
    .X(_3826_));
 sky130_fd_sc_hd__buf_1 _7733_ (.A(_3826_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_2 _7734_ (.A0(_3058_),
    .A1(\rf.registers[30][17] ),
    .S(_3819_),
    .X(_3827_));
 sky130_fd_sc_hd__buf_1 _7735_ (.A(_3827_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_2 _7736_ (.A0(_3060_),
    .A1(\rf.registers[30][18] ),
    .S(_3819_),
    .X(_3828_));
 sky130_fd_sc_hd__buf_1 _7737_ (.A(_3828_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_2 _7738_ (.A0(_3062_),
    .A1(\rf.registers[30][19] ),
    .S(_3819_),
    .X(_3829_));
 sky130_fd_sc_hd__buf_1 _7739_ (.A(_3829_),
    .X(_0361_));
 sky130_fd_sc_hd__buf_1 _7740_ (.A(_3807_),
    .X(_3830_));
 sky130_fd_sc_hd__mux2_2 _7741_ (.A0(_3064_),
    .A1(\rf.registers[30][20] ),
    .S(_3830_),
    .X(_3831_));
 sky130_fd_sc_hd__buf_1 _7742_ (.A(_3831_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_2 _7743_ (.A0(_3067_),
    .A1(\rf.registers[30][21] ),
    .S(_3830_),
    .X(_3832_));
 sky130_fd_sc_hd__buf_1 _7744_ (.A(_3832_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_2 _7745_ (.A0(_3069_),
    .A1(\rf.registers[30][22] ),
    .S(_3830_),
    .X(_3833_));
 sky130_fd_sc_hd__buf_1 _7746_ (.A(_3833_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_2 _7747_ (.A0(_3071_),
    .A1(\rf.registers[30][23] ),
    .S(_3830_),
    .X(_3834_));
 sky130_fd_sc_hd__buf_1 _7748_ (.A(_3834_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_2 _7749_ (.A0(_3073_),
    .A1(\rf.registers[30][24] ),
    .S(_3830_),
    .X(_3835_));
 sky130_fd_sc_hd__buf_1 _7750_ (.A(_3835_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_2 _7751_ (.A0(_3075_),
    .A1(\rf.registers[30][25] ),
    .S(_3830_),
    .X(_3836_));
 sky130_fd_sc_hd__buf_1 _7752_ (.A(_3836_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_2 _7753_ (.A0(_3077_),
    .A1(\rf.registers[30][26] ),
    .S(_3830_),
    .X(_3837_));
 sky130_fd_sc_hd__buf_1 _7754_ (.A(_3837_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_2 _7755_ (.A0(_3079_),
    .A1(\rf.registers[30][27] ),
    .S(_3830_),
    .X(_3838_));
 sky130_fd_sc_hd__buf_1 _7756_ (.A(_3838_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_2 _7757_ (.A0(_3081_),
    .A1(\rf.registers[30][28] ),
    .S(_3830_),
    .X(_3839_));
 sky130_fd_sc_hd__buf_1 _7758_ (.A(_3839_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_2 _7759_ (.A0(_3083_),
    .A1(\rf.registers[30][29] ),
    .S(_3830_),
    .X(_3840_));
 sky130_fd_sc_hd__buf_1 _7760_ (.A(_3840_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_2 _7761_ (.A0(_3085_),
    .A1(\rf.registers[30][30] ),
    .S(_3807_),
    .X(_3841_));
 sky130_fd_sc_hd__buf_1 _7762_ (.A(_3841_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_2 _7763_ (.A0(_3087_),
    .A1(\rf.registers[30][31] ),
    .S(_3807_),
    .X(_3842_));
 sky130_fd_sc_hd__buf_1 _7764_ (.A(_3842_),
    .X(_0373_));
 sky130_fd_sc_hd__nor2_2 _7765_ (.A(_3003_),
    .B(_3091_),
    .Y(_3843_));
 sky130_fd_sc_hd__buf_1 _7766_ (.A(_3843_),
    .X(_3844_));
 sky130_fd_sc_hd__mux2_2 _7767_ (.A0(\rf.registers[9][0] ),
    .A1(_3454_),
    .S(_3844_),
    .X(_3845_));
 sky130_fd_sc_hd__buf_1 _7768_ (.A(_3845_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_2 _7769_ (.A0(\rf.registers[9][1] ),
    .A1(_3458_),
    .S(_3844_),
    .X(_3846_));
 sky130_fd_sc_hd__buf_1 _7770_ (.A(_3846_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_2 _7771_ (.A0(\rf.registers[9][2] ),
    .A1(_3460_),
    .S(_3844_),
    .X(_3847_));
 sky130_fd_sc_hd__buf_1 _7772_ (.A(_3847_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_2 _7773_ (.A0(\rf.registers[9][3] ),
    .A1(_3462_),
    .S(_3844_),
    .X(_3848_));
 sky130_fd_sc_hd__buf_1 _7774_ (.A(_3848_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_2 _7775_ (.A0(\rf.registers[9][4] ),
    .A1(_3464_),
    .S(_3844_),
    .X(_3849_));
 sky130_fd_sc_hd__buf_1 _7776_ (.A(_3849_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_2 _7777_ (.A0(\rf.registers[9][5] ),
    .A1(_3466_),
    .S(_3844_),
    .X(_3850_));
 sky130_fd_sc_hd__buf_1 _7778_ (.A(_3850_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_2 _7779_ (.A0(\rf.registers[9][6] ),
    .A1(_3468_),
    .S(_3844_),
    .X(_3851_));
 sky130_fd_sc_hd__buf_1 _7780_ (.A(_3851_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_2 _7781_ (.A0(\rf.registers[9][7] ),
    .A1(_3470_),
    .S(_3844_),
    .X(_3852_));
 sky130_fd_sc_hd__buf_1 _7782_ (.A(_3852_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_2 _7783_ (.A0(\rf.registers[9][8] ),
    .A1(_3472_),
    .S(_3844_),
    .X(_3853_));
 sky130_fd_sc_hd__buf_1 _7784_ (.A(_3853_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_2 _7785_ (.A0(\rf.registers[9][9] ),
    .A1(_3474_),
    .S(_3844_),
    .X(_3854_));
 sky130_fd_sc_hd__buf_1 _7786_ (.A(_3854_),
    .X(_0383_));
 sky130_fd_sc_hd__buf_1 _7787_ (.A(_3843_),
    .X(_3855_));
 sky130_fd_sc_hd__mux2_2 _7788_ (.A0(\rf.registers[9][10] ),
    .A1(_3476_),
    .S(_3855_),
    .X(_3856_));
 sky130_fd_sc_hd__buf_1 _7789_ (.A(_3856_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_2 _7790_ (.A0(\rf.registers[9][11] ),
    .A1(_3479_),
    .S(_3855_),
    .X(_3857_));
 sky130_fd_sc_hd__buf_1 _7791_ (.A(_3857_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_2 _7792_ (.A0(\rf.registers[9][12] ),
    .A1(_3481_),
    .S(_3855_),
    .X(_3858_));
 sky130_fd_sc_hd__buf_1 _7793_ (.A(_3858_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_2 _7794_ (.A0(\rf.registers[9][13] ),
    .A1(_3483_),
    .S(_3855_),
    .X(_3859_));
 sky130_fd_sc_hd__buf_1 _7795_ (.A(_3859_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_2 _7796_ (.A0(\rf.registers[9][14] ),
    .A1(_3485_),
    .S(_3855_),
    .X(_3860_));
 sky130_fd_sc_hd__buf_1 _7797_ (.A(_3860_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_2 _7798_ (.A0(\rf.registers[9][15] ),
    .A1(_3487_),
    .S(_3855_),
    .X(_3861_));
 sky130_fd_sc_hd__buf_1 _7799_ (.A(_3861_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_2 _7800_ (.A0(\rf.registers[9][16] ),
    .A1(_3489_),
    .S(_3855_),
    .X(_3862_));
 sky130_fd_sc_hd__buf_1 _7801_ (.A(_3862_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_2 _7802_ (.A0(\rf.registers[9][17] ),
    .A1(_3491_),
    .S(_3855_),
    .X(_3863_));
 sky130_fd_sc_hd__buf_1 _7803_ (.A(_3863_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_2 _7804_ (.A0(\rf.registers[9][18] ),
    .A1(_3493_),
    .S(_3855_),
    .X(_3864_));
 sky130_fd_sc_hd__buf_1 _7805_ (.A(_3864_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_2 _7806_ (.A0(\rf.registers[9][19] ),
    .A1(_3495_),
    .S(_3855_),
    .X(_3865_));
 sky130_fd_sc_hd__buf_1 _7807_ (.A(_3865_),
    .X(_0393_));
 sky130_fd_sc_hd__buf_1 _7808_ (.A(_3843_),
    .X(_3866_));
 sky130_fd_sc_hd__mux2_2 _7809_ (.A0(\rf.registers[9][20] ),
    .A1(_3497_),
    .S(_3866_),
    .X(_3867_));
 sky130_fd_sc_hd__buf_1 _7810_ (.A(_3867_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_2 _7811_ (.A0(\rf.registers[9][21] ),
    .A1(_3500_),
    .S(_3866_),
    .X(_3868_));
 sky130_fd_sc_hd__buf_1 _7812_ (.A(_3868_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_2 _7813_ (.A0(\rf.registers[9][22] ),
    .A1(_3502_),
    .S(_3866_),
    .X(_3869_));
 sky130_fd_sc_hd__buf_1 _7814_ (.A(_3869_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_2 _7815_ (.A0(\rf.registers[9][23] ),
    .A1(_3504_),
    .S(_3866_),
    .X(_3870_));
 sky130_fd_sc_hd__buf_1 _7816_ (.A(_3870_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_2 _7817_ (.A0(\rf.registers[9][24] ),
    .A1(_3506_),
    .S(_3866_),
    .X(_3871_));
 sky130_fd_sc_hd__buf_1 _7818_ (.A(_3871_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_2 _7819_ (.A0(\rf.registers[9][25] ),
    .A1(_3508_),
    .S(_3866_),
    .X(_3872_));
 sky130_fd_sc_hd__buf_1 _7820_ (.A(_3872_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_2 _7821_ (.A0(\rf.registers[9][26] ),
    .A1(_3442_),
    .S(_3866_),
    .X(_3873_));
 sky130_fd_sc_hd__buf_1 _7822_ (.A(_3873_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_2 _7823_ (.A0(\rf.registers[9][27] ),
    .A1(_3444_),
    .S(_3866_),
    .X(_3874_));
 sky130_fd_sc_hd__buf_1 _7824_ (.A(_3874_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_2 _7825_ (.A0(\rf.registers[9][28] ),
    .A1(_3446_),
    .S(_3866_),
    .X(_3875_));
 sky130_fd_sc_hd__buf_1 _7826_ (.A(_3875_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_2 _7827_ (.A0(\rf.registers[9][29] ),
    .A1(_3448_),
    .S(_3866_),
    .X(_3876_));
 sky130_fd_sc_hd__buf_1 _7828_ (.A(_3876_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_2 _7829_ (.A0(\rf.registers[9][30] ),
    .A1(_3450_),
    .S(_3843_),
    .X(_3877_));
 sky130_fd_sc_hd__buf_1 _7830_ (.A(_3877_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_2 _7831_ (.A0(\rf.registers[9][31] ),
    .A1(_3452_),
    .S(_3843_),
    .X(_3878_));
 sky130_fd_sc_hd__buf_1 _7832_ (.A(_3878_),
    .X(_0405_));
 sky130_fd_sc_hd__nand2_2 _7833_ (.A(_3021_),
    .B(_3193_),
    .Y(_3879_));
 sky130_fd_sc_hd__buf_1 _7834_ (.A(_3879_),
    .X(_3880_));
 sky130_fd_sc_hd__mux2_2 _7835_ (.A0(_3089_),
    .A1(\rf.registers[23][0] ),
    .S(_3880_),
    .X(_3881_));
 sky130_fd_sc_hd__buf_1 _7836_ (.A(_3881_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_2 _7837_ (.A0(_3095_),
    .A1(\rf.registers[23][1] ),
    .S(_3880_),
    .X(_3882_));
 sky130_fd_sc_hd__buf_1 _7838_ (.A(_3882_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_2 _7839_ (.A0(_3097_),
    .A1(\rf.registers[23][2] ),
    .S(_3880_),
    .X(_3883_));
 sky130_fd_sc_hd__buf_1 _7840_ (.A(_3883_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_2 _7841_ (.A0(_3099_),
    .A1(\rf.registers[23][3] ),
    .S(_3880_),
    .X(_3884_));
 sky130_fd_sc_hd__buf_1 _7842_ (.A(_3884_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_2 _7843_ (.A0(_3101_),
    .A1(\rf.registers[23][4] ),
    .S(_3880_),
    .X(_3885_));
 sky130_fd_sc_hd__buf_1 _7844_ (.A(_3885_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_2 _7845_ (.A0(_3103_),
    .A1(\rf.registers[23][5] ),
    .S(_3880_),
    .X(_3886_));
 sky130_fd_sc_hd__buf_1 _7846_ (.A(_3886_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_2 _7847_ (.A0(_3105_),
    .A1(\rf.registers[23][6] ),
    .S(_3880_),
    .X(_3887_));
 sky130_fd_sc_hd__buf_1 _7848_ (.A(_3887_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_2 _7849_ (.A0(_3107_),
    .A1(\rf.registers[23][7] ),
    .S(_3880_),
    .X(_3888_));
 sky130_fd_sc_hd__buf_1 _7850_ (.A(_3888_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_2 _7851_ (.A0(_3109_),
    .A1(\rf.registers[23][8] ),
    .S(_3880_),
    .X(_3889_));
 sky130_fd_sc_hd__buf_1 _7852_ (.A(_3889_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_2 _7853_ (.A0(_3111_),
    .A1(\rf.registers[23][9] ),
    .S(_3880_),
    .X(_3890_));
 sky130_fd_sc_hd__buf_1 _7854_ (.A(_3890_),
    .X(_0415_));
 sky130_fd_sc_hd__buf_1 _7855_ (.A(_3879_),
    .X(_3891_));
 sky130_fd_sc_hd__mux2_2 _7856_ (.A0(_3113_),
    .A1(\rf.registers[23][10] ),
    .S(_3891_),
    .X(_3892_));
 sky130_fd_sc_hd__buf_1 _7857_ (.A(_3892_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_2 _7858_ (.A0(_3116_),
    .A1(\rf.registers[23][11] ),
    .S(_3891_),
    .X(_3893_));
 sky130_fd_sc_hd__buf_1 _7859_ (.A(_3893_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_2 _7860_ (.A0(_3118_),
    .A1(\rf.registers[23][12] ),
    .S(_3891_),
    .X(_3894_));
 sky130_fd_sc_hd__buf_1 _7861_ (.A(_3894_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_2 _7862_ (.A0(_3120_),
    .A1(\rf.registers[23][13] ),
    .S(_3891_),
    .X(_3895_));
 sky130_fd_sc_hd__buf_1 _7863_ (.A(_3895_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_2 _7864_ (.A0(_3122_),
    .A1(\rf.registers[23][14] ),
    .S(_3891_),
    .X(_3896_));
 sky130_fd_sc_hd__buf_1 _7865_ (.A(_3896_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_2 _7866_ (.A0(_3124_),
    .A1(\rf.registers[23][15] ),
    .S(_3891_),
    .X(_3897_));
 sky130_fd_sc_hd__buf_1 _7867_ (.A(_3897_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_2 _7868_ (.A0(_3126_),
    .A1(\rf.registers[23][16] ),
    .S(_3891_),
    .X(_3898_));
 sky130_fd_sc_hd__buf_1 _7869_ (.A(_3898_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_2 _7870_ (.A0(_3128_),
    .A1(\rf.registers[23][17] ),
    .S(_3891_),
    .X(_3899_));
 sky130_fd_sc_hd__buf_1 _7871_ (.A(_3899_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_2 _7872_ (.A0(_3130_),
    .A1(\rf.registers[23][18] ),
    .S(_3891_),
    .X(_3900_));
 sky130_fd_sc_hd__buf_1 _7873_ (.A(_3900_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_2 _7874_ (.A0(_3132_),
    .A1(\rf.registers[23][19] ),
    .S(_3891_),
    .X(_3901_));
 sky130_fd_sc_hd__buf_1 _7875_ (.A(_3901_),
    .X(_0425_));
 sky130_fd_sc_hd__buf_1 _7876_ (.A(_3879_),
    .X(_3902_));
 sky130_fd_sc_hd__mux2_2 _7877_ (.A0(_3134_),
    .A1(\rf.registers[23][20] ),
    .S(_3902_),
    .X(_3903_));
 sky130_fd_sc_hd__buf_1 _7878_ (.A(_3903_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_2 _7879_ (.A0(_3137_),
    .A1(\rf.registers[23][21] ),
    .S(_3902_),
    .X(_3904_));
 sky130_fd_sc_hd__buf_1 _7880_ (.A(_3904_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_2 _7881_ (.A0(_3139_),
    .A1(\rf.registers[23][22] ),
    .S(_3902_),
    .X(_3905_));
 sky130_fd_sc_hd__buf_1 _7882_ (.A(_3905_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_2 _7883_ (.A0(_3141_),
    .A1(\rf.registers[23][23] ),
    .S(_3902_),
    .X(_3906_));
 sky130_fd_sc_hd__buf_1 _7884_ (.A(_3906_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_2 _7885_ (.A0(_3143_),
    .A1(\rf.registers[23][24] ),
    .S(_3902_),
    .X(_3907_));
 sky130_fd_sc_hd__buf_1 _7886_ (.A(_3907_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_2 _7887_ (.A0(_3145_),
    .A1(\rf.registers[23][25] ),
    .S(_3902_),
    .X(_3908_));
 sky130_fd_sc_hd__buf_1 _7888_ (.A(_3908_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_2 _7889_ (.A0(_3002_),
    .A1(\rf.registers[23][26] ),
    .S(_3902_),
    .X(_3909_));
 sky130_fd_sc_hd__buf_1 _7890_ (.A(_3909_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_2 _7891_ (.A0(_3009_),
    .A1(\rf.registers[23][27] ),
    .S(_3902_),
    .X(_3910_));
 sky130_fd_sc_hd__buf_1 _7892_ (.A(_3910_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_2 _7893_ (.A0(_3011_),
    .A1(\rf.registers[23][28] ),
    .S(_3902_),
    .X(_3911_));
 sky130_fd_sc_hd__buf_1 _7894_ (.A(_3911_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_2 _7895_ (.A0(_3013_),
    .A1(\rf.registers[23][29] ),
    .S(_3902_),
    .X(_3912_));
 sky130_fd_sc_hd__buf_1 _7896_ (.A(_3912_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_2 _7897_ (.A0(_3015_),
    .A1(\rf.registers[23][30] ),
    .S(_3879_),
    .X(_3913_));
 sky130_fd_sc_hd__buf_1 _7898_ (.A(_3913_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_2 _7899_ (.A0(_3017_),
    .A1(\rf.registers[23][31] ),
    .S(_3879_),
    .X(_3914_));
 sky130_fd_sc_hd__buf_1 _7900_ (.A(_3914_),
    .X(_0437_));
 sky130_fd_sc_hd__nor2_2 _7901_ (.A(_3005_),
    .B(_3090_),
    .Y(_3915_));
 sky130_fd_sc_hd__buf_1 _7902_ (.A(_3915_),
    .X(_3916_));
 sky130_fd_sc_hd__mux2_2 _7903_ (.A0(\rf.registers[18][0] ),
    .A1(_3454_),
    .S(_3916_),
    .X(_3917_));
 sky130_fd_sc_hd__buf_1 _7904_ (.A(_3917_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_2 _7905_ (.A0(\rf.registers[18][1] ),
    .A1(_3458_),
    .S(_3916_),
    .X(_3918_));
 sky130_fd_sc_hd__buf_1 _7906_ (.A(_3918_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_2 _7907_ (.A0(\rf.registers[18][2] ),
    .A1(_3460_),
    .S(_3916_),
    .X(_3919_));
 sky130_fd_sc_hd__buf_1 _7908_ (.A(_3919_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_2 _7909_ (.A0(\rf.registers[18][3] ),
    .A1(_3462_),
    .S(_3916_),
    .X(_3920_));
 sky130_fd_sc_hd__buf_1 _7910_ (.A(_3920_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_2 _7911_ (.A0(\rf.registers[18][4] ),
    .A1(_3464_),
    .S(_3916_),
    .X(_3921_));
 sky130_fd_sc_hd__buf_1 _7912_ (.A(_3921_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_2 _7913_ (.A0(\rf.registers[18][5] ),
    .A1(_3466_),
    .S(_3916_),
    .X(_3922_));
 sky130_fd_sc_hd__buf_1 _7914_ (.A(_3922_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_2 _7915_ (.A0(\rf.registers[18][6] ),
    .A1(_3468_),
    .S(_3916_),
    .X(_3923_));
 sky130_fd_sc_hd__buf_1 _7916_ (.A(_3923_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_2 _7917_ (.A0(\rf.registers[18][7] ),
    .A1(_3470_),
    .S(_3916_),
    .X(_3924_));
 sky130_fd_sc_hd__buf_1 _7918_ (.A(_3924_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_2 _7919_ (.A0(\rf.registers[18][8] ),
    .A1(_3472_),
    .S(_3916_),
    .X(_3925_));
 sky130_fd_sc_hd__buf_1 _7920_ (.A(_3925_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_2 _7921_ (.A0(\rf.registers[18][9] ),
    .A1(_3474_),
    .S(_3916_),
    .X(_3926_));
 sky130_fd_sc_hd__buf_1 _7922_ (.A(_3926_),
    .X(_0447_));
 sky130_fd_sc_hd__buf_1 _7923_ (.A(_3915_),
    .X(_3927_));
 sky130_fd_sc_hd__mux2_2 _7924_ (.A0(\rf.registers[18][10] ),
    .A1(_3476_),
    .S(_3927_),
    .X(_3928_));
 sky130_fd_sc_hd__buf_1 _7925_ (.A(_3928_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_2 _7926_ (.A0(\rf.registers[18][11] ),
    .A1(_3479_),
    .S(_3927_),
    .X(_3929_));
 sky130_fd_sc_hd__buf_1 _7927_ (.A(_3929_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_2 _7928_ (.A0(\rf.registers[18][12] ),
    .A1(_3481_),
    .S(_3927_),
    .X(_3930_));
 sky130_fd_sc_hd__buf_1 _7929_ (.A(_3930_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_2 _7930_ (.A0(\rf.registers[18][13] ),
    .A1(_3483_),
    .S(_3927_),
    .X(_3931_));
 sky130_fd_sc_hd__buf_1 _7931_ (.A(_3931_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_2 _7932_ (.A0(\rf.registers[18][14] ),
    .A1(_3485_),
    .S(_3927_),
    .X(_3932_));
 sky130_fd_sc_hd__buf_1 _7933_ (.A(_3932_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_2 _7934_ (.A0(\rf.registers[18][15] ),
    .A1(_3487_),
    .S(_3927_),
    .X(_3933_));
 sky130_fd_sc_hd__buf_1 _7935_ (.A(_3933_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_2 _7936_ (.A0(\rf.registers[18][16] ),
    .A1(_3489_),
    .S(_3927_),
    .X(_3934_));
 sky130_fd_sc_hd__buf_1 _7937_ (.A(_3934_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_2 _7938_ (.A0(\rf.registers[18][17] ),
    .A1(_3491_),
    .S(_3927_),
    .X(_3935_));
 sky130_fd_sc_hd__buf_1 _7939_ (.A(_3935_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_2 _7940_ (.A0(\rf.registers[18][18] ),
    .A1(_3493_),
    .S(_3927_),
    .X(_3936_));
 sky130_fd_sc_hd__buf_1 _7941_ (.A(_3936_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_2 _7942_ (.A0(\rf.registers[18][19] ),
    .A1(_3495_),
    .S(_3927_),
    .X(_3937_));
 sky130_fd_sc_hd__buf_1 _7943_ (.A(_3937_),
    .X(_0457_));
 sky130_fd_sc_hd__buf_1 _7944_ (.A(_3915_),
    .X(_3938_));
 sky130_fd_sc_hd__mux2_2 _7945_ (.A0(\rf.registers[18][20] ),
    .A1(_3497_),
    .S(_3938_),
    .X(_3939_));
 sky130_fd_sc_hd__buf_1 _7946_ (.A(_3939_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_2 _7947_ (.A0(\rf.registers[18][21] ),
    .A1(_3500_),
    .S(_3938_),
    .X(_3940_));
 sky130_fd_sc_hd__buf_1 _7948_ (.A(_3940_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_2 _7949_ (.A0(\rf.registers[18][22] ),
    .A1(_3502_),
    .S(_3938_),
    .X(_3941_));
 sky130_fd_sc_hd__buf_1 _7950_ (.A(_3941_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_2 _7951_ (.A0(\rf.registers[18][23] ),
    .A1(_3504_),
    .S(_3938_),
    .X(_3942_));
 sky130_fd_sc_hd__buf_1 _7952_ (.A(_3942_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_2 _7953_ (.A0(\rf.registers[18][24] ),
    .A1(_3506_),
    .S(_3938_),
    .X(_3943_));
 sky130_fd_sc_hd__buf_1 _7954_ (.A(_3943_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_2 _7955_ (.A0(\rf.registers[18][25] ),
    .A1(_3508_),
    .S(_3938_),
    .X(_3944_));
 sky130_fd_sc_hd__buf_1 _7956_ (.A(_3944_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_2 _7957_ (.A0(\rf.registers[18][26] ),
    .A1(_3442_),
    .S(_3938_),
    .X(_3945_));
 sky130_fd_sc_hd__buf_1 _7958_ (.A(_3945_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_2 _7959_ (.A0(\rf.registers[18][27] ),
    .A1(_3444_),
    .S(_3938_),
    .X(_3946_));
 sky130_fd_sc_hd__buf_1 _7960_ (.A(_3946_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_2 _7961_ (.A0(\rf.registers[18][28] ),
    .A1(_3446_),
    .S(_3938_),
    .X(_3947_));
 sky130_fd_sc_hd__buf_1 _7962_ (.A(_3947_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_2 _7963_ (.A0(\rf.registers[18][29] ),
    .A1(_3448_),
    .S(_3938_),
    .X(_3948_));
 sky130_fd_sc_hd__buf_1 _7964_ (.A(_3948_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_2 _7965_ (.A0(\rf.registers[18][30] ),
    .A1(_3450_),
    .S(_3915_),
    .X(_3949_));
 sky130_fd_sc_hd__buf_1 _7966_ (.A(_3949_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_2 _7967_ (.A0(\rf.registers[18][31] ),
    .A1(_3452_),
    .S(_3915_),
    .X(_3950_));
 sky130_fd_sc_hd__buf_1 _7968_ (.A(_3950_),
    .X(_0469_));
 sky130_fd_sc_hd__nand2_2 _7969_ (.A(_3021_),
    .B(_3552_),
    .Y(_3951_));
 sky130_fd_sc_hd__buf_1 _7970_ (.A(_3951_),
    .X(_3952_));
 sky130_fd_sc_hd__mux2_2 _7971_ (.A0(_3089_),
    .A1(\rf.registers[21][0] ),
    .S(_3952_),
    .X(_3953_));
 sky130_fd_sc_hd__buf_1 _7972_ (.A(_3953_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_2 _7973_ (.A0(_3095_),
    .A1(\rf.registers[21][1] ),
    .S(_3952_),
    .X(_3954_));
 sky130_fd_sc_hd__buf_1 _7974_ (.A(_3954_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_2 _7975_ (.A0(_3097_),
    .A1(\rf.registers[21][2] ),
    .S(_3952_),
    .X(_3955_));
 sky130_fd_sc_hd__buf_1 _7976_ (.A(_3955_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_2 _7977_ (.A0(_3099_),
    .A1(\rf.registers[21][3] ),
    .S(_3952_),
    .X(_3956_));
 sky130_fd_sc_hd__buf_1 _7978_ (.A(_3956_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_2 _7979_ (.A0(_3101_),
    .A1(\rf.registers[21][4] ),
    .S(_3952_),
    .X(_3957_));
 sky130_fd_sc_hd__buf_1 _7980_ (.A(_3957_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_2 _7981_ (.A0(_3103_),
    .A1(\rf.registers[21][5] ),
    .S(_3952_),
    .X(_3958_));
 sky130_fd_sc_hd__buf_1 _7982_ (.A(_3958_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_2 _7983_ (.A0(_3105_),
    .A1(\rf.registers[21][6] ),
    .S(_3952_),
    .X(_3959_));
 sky130_fd_sc_hd__buf_1 _7984_ (.A(_3959_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_2 _7985_ (.A0(_3107_),
    .A1(\rf.registers[21][7] ),
    .S(_3952_),
    .X(_3960_));
 sky130_fd_sc_hd__buf_1 _7986_ (.A(_3960_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_2 _7987_ (.A0(_3109_),
    .A1(\rf.registers[21][8] ),
    .S(_3952_),
    .X(_3961_));
 sky130_fd_sc_hd__buf_1 _7988_ (.A(_3961_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_2 _7989_ (.A0(_3111_),
    .A1(\rf.registers[21][9] ),
    .S(_3952_),
    .X(_3962_));
 sky130_fd_sc_hd__buf_1 _7990_ (.A(_3962_),
    .X(_0479_));
 sky130_fd_sc_hd__buf_1 _7991_ (.A(_3951_),
    .X(_3963_));
 sky130_fd_sc_hd__mux2_2 _7992_ (.A0(_3113_),
    .A1(\rf.registers[21][10] ),
    .S(_3963_),
    .X(_3964_));
 sky130_fd_sc_hd__buf_1 _7993_ (.A(_3964_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_2 _7994_ (.A0(_3116_),
    .A1(\rf.registers[21][11] ),
    .S(_3963_),
    .X(_3965_));
 sky130_fd_sc_hd__buf_1 _7995_ (.A(_3965_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_2 _7996_ (.A0(_3118_),
    .A1(\rf.registers[21][12] ),
    .S(_3963_),
    .X(_3966_));
 sky130_fd_sc_hd__buf_1 _7997_ (.A(_3966_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_2 _7998_ (.A0(_3120_),
    .A1(\rf.registers[21][13] ),
    .S(_3963_),
    .X(_3967_));
 sky130_fd_sc_hd__buf_1 _7999_ (.A(_3967_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_2 _8000_ (.A0(_3122_),
    .A1(\rf.registers[21][14] ),
    .S(_3963_),
    .X(_3968_));
 sky130_fd_sc_hd__buf_1 _8001_ (.A(_3968_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_2 _8002_ (.A0(_3124_),
    .A1(\rf.registers[21][15] ),
    .S(_3963_),
    .X(_3969_));
 sky130_fd_sc_hd__buf_1 _8003_ (.A(_3969_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_2 _8004_ (.A0(_3126_),
    .A1(\rf.registers[21][16] ),
    .S(_3963_),
    .X(_3970_));
 sky130_fd_sc_hd__buf_1 _8005_ (.A(_3970_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_2 _8006_ (.A0(_3128_),
    .A1(\rf.registers[21][17] ),
    .S(_3963_),
    .X(_3971_));
 sky130_fd_sc_hd__buf_1 _8007_ (.A(_3971_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_2 _8008_ (.A0(_3130_),
    .A1(\rf.registers[21][18] ),
    .S(_3963_),
    .X(_3972_));
 sky130_fd_sc_hd__buf_1 _8009_ (.A(_3972_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_2 _8010_ (.A0(_3132_),
    .A1(\rf.registers[21][19] ),
    .S(_3963_),
    .X(_3973_));
 sky130_fd_sc_hd__buf_1 _8011_ (.A(_3973_),
    .X(_0489_));
 sky130_fd_sc_hd__buf_1 _8012_ (.A(_3951_),
    .X(_3974_));
 sky130_fd_sc_hd__mux2_2 _8013_ (.A0(_3134_),
    .A1(\rf.registers[21][20] ),
    .S(_3974_),
    .X(_3975_));
 sky130_fd_sc_hd__buf_1 _8014_ (.A(_3975_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_2 _8015_ (.A0(_3137_),
    .A1(\rf.registers[21][21] ),
    .S(_3974_),
    .X(_3976_));
 sky130_fd_sc_hd__buf_1 _8016_ (.A(_3976_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_2 _8017_ (.A0(_3139_),
    .A1(\rf.registers[21][22] ),
    .S(_3974_),
    .X(_3977_));
 sky130_fd_sc_hd__buf_1 _8018_ (.A(_3977_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_2 _8019_ (.A0(_3141_),
    .A1(\rf.registers[21][23] ),
    .S(_3974_),
    .X(_3978_));
 sky130_fd_sc_hd__buf_1 _8020_ (.A(_3978_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_2 _8021_ (.A0(_3143_),
    .A1(\rf.registers[21][24] ),
    .S(_3974_),
    .X(_3979_));
 sky130_fd_sc_hd__buf_1 _8022_ (.A(_3979_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_2 _8023_ (.A0(_3145_),
    .A1(\rf.registers[21][25] ),
    .S(_3974_),
    .X(_3980_));
 sky130_fd_sc_hd__buf_1 _8024_ (.A(_3980_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_2 _8025_ (.A0(_3002_),
    .A1(\rf.registers[21][26] ),
    .S(_3974_),
    .X(_3981_));
 sky130_fd_sc_hd__buf_1 _8026_ (.A(_3981_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_2 _8027_ (.A0(_3009_),
    .A1(\rf.registers[21][27] ),
    .S(_3974_),
    .X(_3982_));
 sky130_fd_sc_hd__buf_1 _8028_ (.A(_3982_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_2 _8029_ (.A0(_3011_),
    .A1(\rf.registers[21][28] ),
    .S(_3974_),
    .X(_3983_));
 sky130_fd_sc_hd__buf_1 _8030_ (.A(_3983_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_2 _8031_ (.A0(_3013_),
    .A1(\rf.registers[21][29] ),
    .S(_3974_),
    .X(_3984_));
 sky130_fd_sc_hd__buf_1 _8032_ (.A(_3984_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_2 _8033_ (.A0(_3015_),
    .A1(\rf.registers[21][30] ),
    .S(_3951_),
    .X(_3985_));
 sky130_fd_sc_hd__buf_1 _8034_ (.A(_3985_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_2 _8035_ (.A0(_3017_),
    .A1(\rf.registers[21][31] ),
    .S(_3951_),
    .X(_3986_));
 sky130_fd_sc_hd__buf_1 _8036_ (.A(_3986_),
    .X(_0501_));
 sky130_fd_sc_hd__inv_2 _8037_ (.A(_3021_),
    .Y(_3987_));
 sky130_fd_sc_hd__nor2_2 _8038_ (.A(_3987_),
    .B(_3155_),
    .Y(_3988_));
 sky130_fd_sc_hd__buf_1 _8039_ (.A(_3988_),
    .X(_3989_));
 sky130_fd_sc_hd__mux2_2 _8040_ (.A0(\rf.registers[20][0] ),
    .A1(_3454_),
    .S(_3989_),
    .X(_3990_));
 sky130_fd_sc_hd__buf_1 _8041_ (.A(_3990_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_2 _8042_ (.A0(\rf.registers[20][1] ),
    .A1(_3458_),
    .S(_3989_),
    .X(_3991_));
 sky130_fd_sc_hd__buf_1 _8043_ (.A(_3991_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_2 _8044_ (.A0(\rf.registers[20][2] ),
    .A1(_3460_),
    .S(_3989_),
    .X(_3992_));
 sky130_fd_sc_hd__buf_1 _8045_ (.A(_3992_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_2 _8046_ (.A0(\rf.registers[20][3] ),
    .A1(_3462_),
    .S(_3989_),
    .X(_3993_));
 sky130_fd_sc_hd__buf_1 _8047_ (.A(_3993_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_2 _8048_ (.A0(\rf.registers[20][4] ),
    .A1(_3464_),
    .S(_3989_),
    .X(_3994_));
 sky130_fd_sc_hd__buf_1 _8049_ (.A(_3994_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_2 _8050_ (.A0(\rf.registers[20][5] ),
    .A1(_3466_),
    .S(_3989_),
    .X(_3995_));
 sky130_fd_sc_hd__buf_1 _8051_ (.A(_3995_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_2 _8052_ (.A0(\rf.registers[20][6] ),
    .A1(_3468_),
    .S(_3989_),
    .X(_3996_));
 sky130_fd_sc_hd__buf_1 _8053_ (.A(_3996_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_2 _8054_ (.A0(\rf.registers[20][7] ),
    .A1(_3470_),
    .S(_3989_),
    .X(_3997_));
 sky130_fd_sc_hd__buf_1 _8055_ (.A(_3997_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_2 _8056_ (.A0(\rf.registers[20][8] ),
    .A1(_3472_),
    .S(_3989_),
    .X(_3998_));
 sky130_fd_sc_hd__buf_1 _8057_ (.A(_3998_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_2 _8058_ (.A0(\rf.registers[20][9] ),
    .A1(_3474_),
    .S(_3989_),
    .X(_3999_));
 sky130_fd_sc_hd__buf_1 _8059_ (.A(_3999_),
    .X(_0511_));
 sky130_fd_sc_hd__buf_1 _8060_ (.A(_3988_),
    .X(_4000_));
 sky130_fd_sc_hd__mux2_2 _8061_ (.A0(\rf.registers[20][10] ),
    .A1(_3476_),
    .S(_4000_),
    .X(_4001_));
 sky130_fd_sc_hd__buf_1 _8062_ (.A(_4001_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_2 _8063_ (.A0(\rf.registers[20][11] ),
    .A1(_3479_),
    .S(_4000_),
    .X(_4002_));
 sky130_fd_sc_hd__buf_1 _8064_ (.A(_4002_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_2 _8065_ (.A0(\rf.registers[20][12] ),
    .A1(_3481_),
    .S(_4000_),
    .X(_4003_));
 sky130_fd_sc_hd__buf_1 _8066_ (.A(_4003_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_2 _8067_ (.A0(\rf.registers[20][13] ),
    .A1(_3483_),
    .S(_4000_),
    .X(_4004_));
 sky130_fd_sc_hd__buf_1 _8068_ (.A(_4004_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_2 _8069_ (.A0(\rf.registers[20][14] ),
    .A1(_3485_),
    .S(_4000_),
    .X(_4005_));
 sky130_fd_sc_hd__buf_1 _8070_ (.A(_4005_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_2 _8071_ (.A0(\rf.registers[20][15] ),
    .A1(_3487_),
    .S(_4000_),
    .X(_4006_));
 sky130_fd_sc_hd__buf_1 _8072_ (.A(_4006_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_2 _8073_ (.A0(\rf.registers[20][16] ),
    .A1(_3489_),
    .S(_4000_),
    .X(_4007_));
 sky130_fd_sc_hd__buf_1 _8074_ (.A(_4007_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_2 _8075_ (.A0(\rf.registers[20][17] ),
    .A1(_3491_),
    .S(_4000_),
    .X(_4008_));
 sky130_fd_sc_hd__buf_1 _8076_ (.A(_4008_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_2 _8077_ (.A0(\rf.registers[20][18] ),
    .A1(_3493_),
    .S(_4000_),
    .X(_4009_));
 sky130_fd_sc_hd__buf_1 _8078_ (.A(_4009_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_2 _8079_ (.A0(\rf.registers[20][19] ),
    .A1(_3495_),
    .S(_4000_),
    .X(_4010_));
 sky130_fd_sc_hd__buf_1 _8080_ (.A(_4010_),
    .X(_0521_));
 sky130_fd_sc_hd__buf_1 _8081_ (.A(_3988_),
    .X(_4011_));
 sky130_fd_sc_hd__mux2_2 _8082_ (.A0(\rf.registers[20][20] ),
    .A1(_3497_),
    .S(_4011_),
    .X(_4012_));
 sky130_fd_sc_hd__buf_1 _8083_ (.A(_4012_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_2 _8084_ (.A0(\rf.registers[20][21] ),
    .A1(_3500_),
    .S(_4011_),
    .X(_4013_));
 sky130_fd_sc_hd__buf_1 _8085_ (.A(_4013_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_2 _8086_ (.A0(\rf.registers[20][22] ),
    .A1(_3502_),
    .S(_4011_),
    .X(_4014_));
 sky130_fd_sc_hd__buf_1 _8087_ (.A(_4014_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_2 _8088_ (.A0(\rf.registers[20][23] ),
    .A1(_3504_),
    .S(_4011_),
    .X(_4015_));
 sky130_fd_sc_hd__buf_1 _8089_ (.A(_4015_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_2 _8090_ (.A0(\rf.registers[20][24] ),
    .A1(_3506_),
    .S(_4011_),
    .X(_4016_));
 sky130_fd_sc_hd__buf_1 _8091_ (.A(_4016_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_2 _8092_ (.A0(\rf.registers[20][25] ),
    .A1(_3508_),
    .S(_4011_),
    .X(_4017_));
 sky130_fd_sc_hd__buf_1 _8093_ (.A(_4017_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_2 _8094_ (.A0(\rf.registers[20][26] ),
    .A1(_3442_),
    .S(_4011_),
    .X(_4018_));
 sky130_fd_sc_hd__buf_1 _8095_ (.A(_4018_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_2 _8096_ (.A0(\rf.registers[20][27] ),
    .A1(_3444_),
    .S(_4011_),
    .X(_4019_));
 sky130_fd_sc_hd__buf_1 _8097_ (.A(_4019_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_2 _8098_ (.A0(\rf.registers[20][28] ),
    .A1(_3446_),
    .S(_4011_),
    .X(_4020_));
 sky130_fd_sc_hd__buf_1 _8099_ (.A(_4020_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_2 _8100_ (.A0(\rf.registers[20][29] ),
    .A1(_3448_),
    .S(_4011_),
    .X(_4021_));
 sky130_fd_sc_hd__buf_1 _8101_ (.A(_4021_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_2 _8102_ (.A0(\rf.registers[20][30] ),
    .A1(_3450_),
    .S(_3988_),
    .X(_4022_));
 sky130_fd_sc_hd__buf_1 _8103_ (.A(_4022_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_2 _8104_ (.A0(\rf.registers[20][31] ),
    .A1(_3452_),
    .S(_3988_),
    .X(_4023_));
 sky130_fd_sc_hd__buf_1 _8105_ (.A(_4023_),
    .X(_0533_));
 sky130_fd_sc_hd__nor2b_2 _8106_ (.A(_3155_),
    .B_N(_3626_),
    .Y(_4024_));
 sky130_fd_sc_hd__buf_1 _8107_ (.A(_4024_),
    .X(_4025_));
 sky130_fd_sc_hd__mux2_2 _8108_ (.A0(\rf.registers[24][0] ),
    .A1(_3454_),
    .S(_4025_),
    .X(_4026_));
 sky130_fd_sc_hd__buf_1 _8109_ (.A(_4026_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_2 _8110_ (.A0(\rf.registers[24][1] ),
    .A1(_3458_),
    .S(_4025_),
    .X(_4027_));
 sky130_fd_sc_hd__buf_1 _8111_ (.A(_4027_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_2 _8112_ (.A0(\rf.registers[24][2] ),
    .A1(_3460_),
    .S(_4025_),
    .X(_4028_));
 sky130_fd_sc_hd__buf_1 _8113_ (.A(_4028_),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_2 _8114_ (.A0(\rf.registers[24][3] ),
    .A1(_3462_),
    .S(_4025_),
    .X(_4029_));
 sky130_fd_sc_hd__buf_1 _8115_ (.A(_4029_),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_2 _8116_ (.A0(\rf.registers[24][4] ),
    .A1(_3464_),
    .S(_4025_),
    .X(_4030_));
 sky130_fd_sc_hd__buf_1 _8117_ (.A(_4030_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_2 _8118_ (.A0(\rf.registers[24][5] ),
    .A1(_3466_),
    .S(_4025_),
    .X(_4031_));
 sky130_fd_sc_hd__buf_1 _8119_ (.A(_4031_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_2 _8120_ (.A0(\rf.registers[24][6] ),
    .A1(_3468_),
    .S(_4025_),
    .X(_4032_));
 sky130_fd_sc_hd__buf_1 _8121_ (.A(_4032_),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_2 _8122_ (.A0(\rf.registers[24][7] ),
    .A1(_3470_),
    .S(_4025_),
    .X(_4033_));
 sky130_fd_sc_hd__buf_1 _8123_ (.A(_4033_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_2 _8124_ (.A0(\rf.registers[24][8] ),
    .A1(_3472_),
    .S(_4025_),
    .X(_4034_));
 sky130_fd_sc_hd__buf_1 _8125_ (.A(_4034_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_2 _8126_ (.A0(\rf.registers[24][9] ),
    .A1(_3474_),
    .S(_4025_),
    .X(_4035_));
 sky130_fd_sc_hd__buf_1 _8127_ (.A(_4035_),
    .X(_0543_));
 sky130_fd_sc_hd__buf_1 _8128_ (.A(_4024_),
    .X(_4036_));
 sky130_fd_sc_hd__mux2_2 _8129_ (.A0(\rf.registers[24][10] ),
    .A1(_3476_),
    .S(_4036_),
    .X(_4037_));
 sky130_fd_sc_hd__buf_1 _8130_ (.A(_4037_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_2 _8131_ (.A0(\rf.registers[24][11] ),
    .A1(_3479_),
    .S(_4036_),
    .X(_4038_));
 sky130_fd_sc_hd__buf_1 _8132_ (.A(_4038_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_2 _8133_ (.A0(\rf.registers[24][12] ),
    .A1(_3481_),
    .S(_4036_),
    .X(_4039_));
 sky130_fd_sc_hd__buf_1 _8134_ (.A(_4039_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_2 _8135_ (.A0(\rf.registers[24][13] ),
    .A1(_3483_),
    .S(_4036_),
    .X(_4040_));
 sky130_fd_sc_hd__buf_1 _8136_ (.A(_4040_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_2 _8137_ (.A0(\rf.registers[24][14] ),
    .A1(_3485_),
    .S(_4036_),
    .X(_4041_));
 sky130_fd_sc_hd__buf_1 _8138_ (.A(_4041_),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_2 _8139_ (.A0(\rf.registers[24][15] ),
    .A1(_3487_),
    .S(_4036_),
    .X(_4042_));
 sky130_fd_sc_hd__buf_1 _8140_ (.A(_4042_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_2 _8141_ (.A0(\rf.registers[24][16] ),
    .A1(_3489_),
    .S(_4036_),
    .X(_4043_));
 sky130_fd_sc_hd__buf_1 _8142_ (.A(_4043_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_2 _8143_ (.A0(\rf.registers[24][17] ),
    .A1(_3491_),
    .S(_4036_),
    .X(_4044_));
 sky130_fd_sc_hd__buf_1 _8144_ (.A(_4044_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_2 _8145_ (.A0(\rf.registers[24][18] ),
    .A1(_3493_),
    .S(_4036_),
    .X(_4045_));
 sky130_fd_sc_hd__buf_1 _8146_ (.A(_4045_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_2 _8147_ (.A0(\rf.registers[24][19] ),
    .A1(_3495_),
    .S(_4036_),
    .X(_4046_));
 sky130_fd_sc_hd__buf_1 _8148_ (.A(_4046_),
    .X(_0553_));
 sky130_fd_sc_hd__buf_1 _8149_ (.A(_4024_),
    .X(_4047_));
 sky130_fd_sc_hd__mux2_2 _8150_ (.A0(\rf.registers[24][20] ),
    .A1(_3497_),
    .S(_4047_),
    .X(_4048_));
 sky130_fd_sc_hd__buf_1 _8151_ (.A(_4048_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_2 _8152_ (.A0(\rf.registers[24][21] ),
    .A1(_3500_),
    .S(_4047_),
    .X(_4049_));
 sky130_fd_sc_hd__buf_1 _8153_ (.A(_4049_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_2 _8154_ (.A0(\rf.registers[24][22] ),
    .A1(_3502_),
    .S(_4047_),
    .X(_4050_));
 sky130_fd_sc_hd__buf_1 _8155_ (.A(_4050_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_2 _8156_ (.A0(\rf.registers[24][23] ),
    .A1(_3504_),
    .S(_4047_),
    .X(_4051_));
 sky130_fd_sc_hd__buf_1 _8157_ (.A(_4051_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_2 _8158_ (.A0(\rf.registers[24][24] ),
    .A1(_3506_),
    .S(_4047_),
    .X(_4052_));
 sky130_fd_sc_hd__buf_1 _8159_ (.A(_4052_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_2 _8160_ (.A0(\rf.registers[24][25] ),
    .A1(_3508_),
    .S(_4047_),
    .X(_4053_));
 sky130_fd_sc_hd__buf_1 _8161_ (.A(_4053_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_2 _8162_ (.A0(\rf.registers[24][26] ),
    .A1(_3442_),
    .S(_4047_),
    .X(_4054_));
 sky130_fd_sc_hd__buf_1 _8163_ (.A(_4054_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_2 _8164_ (.A0(\rf.registers[24][27] ),
    .A1(_3444_),
    .S(_4047_),
    .X(_4055_));
 sky130_fd_sc_hd__buf_1 _8165_ (.A(_4055_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_2 _8166_ (.A0(\rf.registers[24][28] ),
    .A1(_3446_),
    .S(_4047_),
    .X(_4056_));
 sky130_fd_sc_hd__buf_1 _8167_ (.A(_4056_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_2 _8168_ (.A0(\rf.registers[24][29] ),
    .A1(_3448_),
    .S(_4047_),
    .X(_4057_));
 sky130_fd_sc_hd__buf_1 _8169_ (.A(_4057_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_2 _8170_ (.A0(\rf.registers[24][30] ),
    .A1(_3450_),
    .S(_4024_),
    .X(_4058_));
 sky130_fd_sc_hd__buf_1 _8171_ (.A(_4058_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_2 _8172_ (.A0(\rf.registers[24][31] ),
    .A1(_3452_),
    .S(_4024_),
    .X(_4059_));
 sky130_fd_sc_hd__buf_1 _8173_ (.A(_4059_),
    .X(_0565_));
 sky130_fd_sc_hd__nor2_2 _8174_ (.A(_3091_),
    .B(_3153_),
    .Y(_4060_));
 sky130_fd_sc_hd__buf_1 _8175_ (.A(_4060_),
    .X(_4061_));
 sky130_fd_sc_hd__mux2_2 _8176_ (.A0(\rf.registers[1][0] ),
    .A1(_3454_),
    .S(_4061_),
    .X(_4062_));
 sky130_fd_sc_hd__buf_1 _8177_ (.A(_4062_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_2 _8178_ (.A0(\rf.registers[1][1] ),
    .A1(_3458_),
    .S(_4061_),
    .X(_4063_));
 sky130_fd_sc_hd__buf_1 _8179_ (.A(_4063_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_2 _8180_ (.A0(\rf.registers[1][2] ),
    .A1(_3460_),
    .S(_4061_),
    .X(_4064_));
 sky130_fd_sc_hd__buf_1 _8181_ (.A(_4064_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_2 _8182_ (.A0(\rf.registers[1][3] ),
    .A1(_3462_),
    .S(_4061_),
    .X(_4065_));
 sky130_fd_sc_hd__buf_1 _8183_ (.A(_4065_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_2 _8184_ (.A0(\rf.registers[1][4] ),
    .A1(_3464_),
    .S(_4061_),
    .X(_4066_));
 sky130_fd_sc_hd__buf_1 _8185_ (.A(_4066_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_2 _8186_ (.A0(\rf.registers[1][5] ),
    .A1(_3466_),
    .S(_4061_),
    .X(_4067_));
 sky130_fd_sc_hd__buf_1 _8187_ (.A(_4067_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_2 _8188_ (.A0(\rf.registers[1][6] ),
    .A1(_3468_),
    .S(_4061_),
    .X(_4068_));
 sky130_fd_sc_hd__buf_1 _8189_ (.A(_4068_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_2 _8190_ (.A0(\rf.registers[1][7] ),
    .A1(_3470_),
    .S(_4061_),
    .X(_4069_));
 sky130_fd_sc_hd__buf_1 _8191_ (.A(_4069_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_2 _8192_ (.A0(\rf.registers[1][8] ),
    .A1(_3472_),
    .S(_4061_),
    .X(_4070_));
 sky130_fd_sc_hd__buf_1 _8193_ (.A(_4070_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_2 _8194_ (.A0(\rf.registers[1][9] ),
    .A1(_3474_),
    .S(_4061_),
    .X(_4071_));
 sky130_fd_sc_hd__buf_1 _8195_ (.A(_4071_),
    .X(_0575_));
 sky130_fd_sc_hd__buf_1 _8196_ (.A(_4060_),
    .X(_4072_));
 sky130_fd_sc_hd__mux2_2 _8197_ (.A0(\rf.registers[1][10] ),
    .A1(_3476_),
    .S(_4072_),
    .X(_4073_));
 sky130_fd_sc_hd__buf_1 _8198_ (.A(_4073_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_2 _8199_ (.A0(\rf.registers[1][11] ),
    .A1(_3479_),
    .S(_4072_),
    .X(_4074_));
 sky130_fd_sc_hd__buf_1 _8200_ (.A(_4074_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_2 _8201_ (.A0(\rf.registers[1][12] ),
    .A1(_3481_),
    .S(_4072_),
    .X(_4075_));
 sky130_fd_sc_hd__buf_1 _8202_ (.A(_4075_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_2 _8203_ (.A0(\rf.registers[1][13] ),
    .A1(_3483_),
    .S(_4072_),
    .X(_4076_));
 sky130_fd_sc_hd__buf_1 _8204_ (.A(_4076_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_2 _8205_ (.A0(\rf.registers[1][14] ),
    .A1(_3485_),
    .S(_4072_),
    .X(_4077_));
 sky130_fd_sc_hd__buf_1 _8206_ (.A(_4077_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_2 _8207_ (.A0(\rf.registers[1][15] ),
    .A1(_3487_),
    .S(_4072_),
    .X(_4078_));
 sky130_fd_sc_hd__buf_1 _8208_ (.A(_4078_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_2 _8209_ (.A0(\rf.registers[1][16] ),
    .A1(_3489_),
    .S(_4072_),
    .X(_4079_));
 sky130_fd_sc_hd__buf_1 _8210_ (.A(_4079_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_2 _8211_ (.A0(\rf.registers[1][17] ),
    .A1(_3491_),
    .S(_4072_),
    .X(_4080_));
 sky130_fd_sc_hd__buf_1 _8212_ (.A(_4080_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_2 _8213_ (.A0(\rf.registers[1][18] ),
    .A1(_3493_),
    .S(_4072_),
    .X(_4081_));
 sky130_fd_sc_hd__buf_1 _8214_ (.A(_4081_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_2 _8215_ (.A0(\rf.registers[1][19] ),
    .A1(_3495_),
    .S(_4072_),
    .X(_4082_));
 sky130_fd_sc_hd__buf_1 _8216_ (.A(_4082_),
    .X(_0585_));
 sky130_fd_sc_hd__buf_1 _8217_ (.A(_4060_),
    .X(_4083_));
 sky130_fd_sc_hd__mux2_2 _8218_ (.A0(\rf.registers[1][20] ),
    .A1(_3497_),
    .S(_4083_),
    .X(_4084_));
 sky130_fd_sc_hd__buf_1 _8219_ (.A(_4084_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_2 _8220_ (.A0(\rf.registers[1][21] ),
    .A1(_3500_),
    .S(_4083_),
    .X(_4085_));
 sky130_fd_sc_hd__buf_1 _8221_ (.A(_4085_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_2 _8222_ (.A0(\rf.registers[1][22] ),
    .A1(_3502_),
    .S(_4083_),
    .X(_4086_));
 sky130_fd_sc_hd__buf_1 _8223_ (.A(_4086_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_2 _8224_ (.A0(\rf.registers[1][23] ),
    .A1(_3504_),
    .S(_4083_),
    .X(_4087_));
 sky130_fd_sc_hd__buf_1 _8225_ (.A(_4087_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_2 _8226_ (.A0(\rf.registers[1][24] ),
    .A1(_3506_),
    .S(_4083_),
    .X(_4088_));
 sky130_fd_sc_hd__buf_1 _8227_ (.A(_4088_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_2 _8228_ (.A0(\rf.registers[1][25] ),
    .A1(_3508_),
    .S(_4083_),
    .X(_4089_));
 sky130_fd_sc_hd__buf_1 _8229_ (.A(_4089_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_2 _8230_ (.A0(\rf.registers[1][26] ),
    .A1(_3442_),
    .S(_4083_),
    .X(_4090_));
 sky130_fd_sc_hd__buf_1 _8231_ (.A(_4090_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_2 _8232_ (.A0(\rf.registers[1][27] ),
    .A1(_3444_),
    .S(_4083_),
    .X(_4091_));
 sky130_fd_sc_hd__buf_1 _8233_ (.A(_4091_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_2 _8234_ (.A0(\rf.registers[1][28] ),
    .A1(_3446_),
    .S(_4083_),
    .X(_4092_));
 sky130_fd_sc_hd__buf_1 _8235_ (.A(_4092_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_2 _8236_ (.A0(\rf.registers[1][29] ),
    .A1(_3448_),
    .S(_4083_),
    .X(_4093_));
 sky130_fd_sc_hd__buf_1 _8237_ (.A(_4093_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_2 _8238_ (.A0(\rf.registers[1][30] ),
    .A1(_3450_),
    .S(_4060_),
    .X(_4094_));
 sky130_fd_sc_hd__buf_1 _8239_ (.A(_4094_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_2 _8240_ (.A0(\rf.registers[1][31] ),
    .A1(_3452_),
    .S(_4060_),
    .X(_4095_));
 sky130_fd_sc_hd__buf_1 _8241_ (.A(_4095_),
    .X(_0597_));
 sky130_fd_sc_hd__nand2_2 _8242_ (.A(_3552_),
    .B(_3192_),
    .Y(_4096_));
 sky130_fd_sc_hd__buf_1 _8243_ (.A(_4096_),
    .X(_4097_));
 sky130_fd_sc_hd__mux2_2 _8244_ (.A0(_3089_),
    .A1(\rf.registers[13][0] ),
    .S(_4097_),
    .X(_4098_));
 sky130_fd_sc_hd__buf_1 _8245_ (.A(_4098_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_2 _8246_ (.A0(_3095_),
    .A1(\rf.registers[13][1] ),
    .S(_4097_),
    .X(_4099_));
 sky130_fd_sc_hd__buf_1 _8247_ (.A(_4099_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_2 _8248_ (.A0(_3097_),
    .A1(\rf.registers[13][2] ),
    .S(_4097_),
    .X(_4100_));
 sky130_fd_sc_hd__buf_1 _8249_ (.A(_4100_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_2 _8250_ (.A0(_3099_),
    .A1(\rf.registers[13][3] ),
    .S(_4097_),
    .X(_4101_));
 sky130_fd_sc_hd__buf_1 _8251_ (.A(_4101_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_2 _8252_ (.A0(_3101_),
    .A1(\rf.registers[13][4] ),
    .S(_4097_),
    .X(_4102_));
 sky130_fd_sc_hd__buf_1 _8253_ (.A(_4102_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_2 _8254_ (.A0(_3103_),
    .A1(\rf.registers[13][5] ),
    .S(_4097_),
    .X(_4103_));
 sky130_fd_sc_hd__buf_1 _8255_ (.A(_4103_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_2 _8256_ (.A0(_3105_),
    .A1(\rf.registers[13][6] ),
    .S(_4097_),
    .X(_4104_));
 sky130_fd_sc_hd__buf_1 _8257_ (.A(_4104_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_2 _8258_ (.A0(_3107_),
    .A1(\rf.registers[13][7] ),
    .S(_4097_),
    .X(_4105_));
 sky130_fd_sc_hd__buf_1 _8259_ (.A(_4105_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_2 _8260_ (.A0(_3109_),
    .A1(\rf.registers[13][8] ),
    .S(_4097_),
    .X(_4106_));
 sky130_fd_sc_hd__buf_1 _8261_ (.A(_4106_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_2 _8262_ (.A0(_3111_),
    .A1(\rf.registers[13][9] ),
    .S(_4097_),
    .X(_4107_));
 sky130_fd_sc_hd__buf_1 _8263_ (.A(_4107_),
    .X(_0607_));
 sky130_fd_sc_hd__buf_1 _8264_ (.A(_4096_),
    .X(_4108_));
 sky130_fd_sc_hd__mux2_2 _8265_ (.A0(_3113_),
    .A1(\rf.registers[13][10] ),
    .S(_4108_),
    .X(_4109_));
 sky130_fd_sc_hd__buf_1 _8266_ (.A(_4109_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_2 _8267_ (.A0(_3116_),
    .A1(\rf.registers[13][11] ),
    .S(_4108_),
    .X(_4110_));
 sky130_fd_sc_hd__buf_1 _8268_ (.A(_4110_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_2 _8269_ (.A0(_3118_),
    .A1(\rf.registers[13][12] ),
    .S(_4108_),
    .X(_4111_));
 sky130_fd_sc_hd__buf_1 _8270_ (.A(_4111_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_2 _8271_ (.A0(_3120_),
    .A1(\rf.registers[13][13] ),
    .S(_4108_),
    .X(_4112_));
 sky130_fd_sc_hd__buf_1 _8272_ (.A(_4112_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_2 _8273_ (.A0(_3122_),
    .A1(\rf.registers[13][14] ),
    .S(_4108_),
    .X(_4113_));
 sky130_fd_sc_hd__buf_1 _8274_ (.A(_4113_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_2 _8275_ (.A0(_3124_),
    .A1(\rf.registers[13][15] ),
    .S(_4108_),
    .X(_4114_));
 sky130_fd_sc_hd__buf_1 _8276_ (.A(_4114_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_2 _8277_ (.A0(_3126_),
    .A1(\rf.registers[13][16] ),
    .S(_4108_),
    .X(_4115_));
 sky130_fd_sc_hd__buf_1 _8278_ (.A(_4115_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_2 _8279_ (.A0(_3128_),
    .A1(\rf.registers[13][17] ),
    .S(_4108_),
    .X(_4116_));
 sky130_fd_sc_hd__buf_1 _8280_ (.A(_4116_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_2 _8281_ (.A0(_3130_),
    .A1(\rf.registers[13][18] ),
    .S(_4108_),
    .X(_4117_));
 sky130_fd_sc_hd__buf_1 _8282_ (.A(_4117_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_2 _8283_ (.A0(_3132_),
    .A1(\rf.registers[13][19] ),
    .S(_4108_),
    .X(_4118_));
 sky130_fd_sc_hd__buf_1 _8284_ (.A(_4118_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_1 _8285_ (.A(_4096_),
    .X(_4119_));
 sky130_fd_sc_hd__mux2_2 _8286_ (.A0(_3134_),
    .A1(\rf.registers[13][20] ),
    .S(_4119_),
    .X(_4120_));
 sky130_fd_sc_hd__buf_1 _8287_ (.A(_4120_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_2 _8288_ (.A0(_3137_),
    .A1(\rf.registers[13][21] ),
    .S(_4119_),
    .X(_4121_));
 sky130_fd_sc_hd__buf_1 _8289_ (.A(_4121_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_2 _8290_ (.A0(_3139_),
    .A1(\rf.registers[13][22] ),
    .S(_4119_),
    .X(_4122_));
 sky130_fd_sc_hd__buf_1 _8291_ (.A(_4122_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_2 _8292_ (.A0(_3141_),
    .A1(\rf.registers[13][23] ),
    .S(_4119_),
    .X(_4123_));
 sky130_fd_sc_hd__buf_1 _8293_ (.A(_4123_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_2 _8294_ (.A0(_3143_),
    .A1(\rf.registers[13][24] ),
    .S(_4119_),
    .X(_4124_));
 sky130_fd_sc_hd__buf_1 _8295_ (.A(_4124_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_2 _8296_ (.A0(_3145_),
    .A1(\rf.registers[13][25] ),
    .S(_4119_),
    .X(_4125_));
 sky130_fd_sc_hd__buf_1 _8297_ (.A(_4125_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_2 _8298_ (.A0(_3002_),
    .A1(\rf.registers[13][26] ),
    .S(_4119_),
    .X(_4126_));
 sky130_fd_sc_hd__buf_1 _8299_ (.A(_4126_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_2 _8300_ (.A0(_3009_),
    .A1(\rf.registers[13][27] ),
    .S(_4119_),
    .X(_4127_));
 sky130_fd_sc_hd__buf_1 _8301_ (.A(_4127_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_2 _8302_ (.A0(_3011_),
    .A1(\rf.registers[13][28] ),
    .S(_4119_),
    .X(_4128_));
 sky130_fd_sc_hd__buf_1 _8303_ (.A(_4128_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_2 _8304_ (.A0(_3013_),
    .A1(\rf.registers[13][29] ),
    .S(_4119_),
    .X(_4129_));
 sky130_fd_sc_hd__buf_1 _8305_ (.A(_4129_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_2 _8306_ (.A0(_3015_),
    .A1(\rf.registers[13][30] ),
    .S(_4096_),
    .X(_4130_));
 sky130_fd_sc_hd__buf_1 _8307_ (.A(_4130_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_2 _8308_ (.A0(_3017_),
    .A1(\rf.registers[13][31] ),
    .S(_4096_),
    .X(_4131_));
 sky130_fd_sc_hd__buf_1 _8309_ (.A(_4131_),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_2 _8310_ (.A(_3090_),
    .B(_3155_),
    .Y(_4132_));
 sky130_fd_sc_hd__buf_1 _8311_ (.A(_4132_),
    .X(_4133_));
 sky130_fd_sc_hd__mux2_2 _8312_ (.A0(\rf.registers[16][0] ),
    .A1(_3454_),
    .S(_4133_),
    .X(_4134_));
 sky130_fd_sc_hd__buf_1 _8313_ (.A(_4134_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_2 _8314_ (.A0(\rf.registers[16][1] ),
    .A1(_3458_),
    .S(_4133_),
    .X(_4135_));
 sky130_fd_sc_hd__buf_1 _8315_ (.A(_4135_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_2 _8316_ (.A0(\rf.registers[16][2] ),
    .A1(_3460_),
    .S(_4133_),
    .X(_4136_));
 sky130_fd_sc_hd__buf_1 _8317_ (.A(_4136_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_2 _8318_ (.A0(\rf.registers[16][3] ),
    .A1(_3462_),
    .S(_4133_),
    .X(_4137_));
 sky130_fd_sc_hd__buf_1 _8319_ (.A(_4137_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_2 _8320_ (.A0(\rf.registers[16][4] ),
    .A1(_3464_),
    .S(_4133_),
    .X(_4138_));
 sky130_fd_sc_hd__buf_1 _8321_ (.A(_4138_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_2 _8322_ (.A0(\rf.registers[16][5] ),
    .A1(_3466_),
    .S(_4133_),
    .X(_4139_));
 sky130_fd_sc_hd__buf_1 _8323_ (.A(_4139_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_2 _8324_ (.A0(\rf.registers[16][6] ),
    .A1(_3468_),
    .S(_4133_),
    .X(_4140_));
 sky130_fd_sc_hd__buf_1 _8325_ (.A(_4140_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_2 _8326_ (.A0(\rf.registers[16][7] ),
    .A1(_3470_),
    .S(_4133_),
    .X(_4141_));
 sky130_fd_sc_hd__buf_1 _8327_ (.A(_4141_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_2 _8328_ (.A0(\rf.registers[16][8] ),
    .A1(_3472_),
    .S(_4133_),
    .X(_4142_));
 sky130_fd_sc_hd__buf_1 _8329_ (.A(_4142_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_2 _8330_ (.A0(\rf.registers[16][9] ),
    .A1(_3474_),
    .S(_4133_),
    .X(_4143_));
 sky130_fd_sc_hd__buf_1 _8331_ (.A(_4143_),
    .X(_0639_));
 sky130_fd_sc_hd__buf_1 _8332_ (.A(_4132_),
    .X(_4144_));
 sky130_fd_sc_hd__mux2_2 _8333_ (.A0(\rf.registers[16][10] ),
    .A1(_3476_),
    .S(_4144_),
    .X(_4145_));
 sky130_fd_sc_hd__buf_1 _8334_ (.A(_4145_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_2 _8335_ (.A0(\rf.registers[16][11] ),
    .A1(_3479_),
    .S(_4144_),
    .X(_4146_));
 sky130_fd_sc_hd__buf_1 _8336_ (.A(_4146_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_2 _8337_ (.A0(\rf.registers[16][12] ),
    .A1(_3481_),
    .S(_4144_),
    .X(_4147_));
 sky130_fd_sc_hd__buf_1 _8338_ (.A(_4147_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_2 _8339_ (.A0(\rf.registers[16][13] ),
    .A1(_3483_),
    .S(_4144_),
    .X(_4148_));
 sky130_fd_sc_hd__buf_1 _8340_ (.A(_4148_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_2 _8341_ (.A0(\rf.registers[16][14] ),
    .A1(_3485_),
    .S(_4144_),
    .X(_4149_));
 sky130_fd_sc_hd__buf_1 _8342_ (.A(_4149_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_2 _8343_ (.A0(\rf.registers[16][15] ),
    .A1(_3487_),
    .S(_4144_),
    .X(_4150_));
 sky130_fd_sc_hd__buf_1 _8344_ (.A(_4150_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_2 _8345_ (.A0(\rf.registers[16][16] ),
    .A1(_3489_),
    .S(_4144_),
    .X(_4151_));
 sky130_fd_sc_hd__buf_1 _8346_ (.A(_4151_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_2 _8347_ (.A0(\rf.registers[16][17] ),
    .A1(_3491_),
    .S(_4144_),
    .X(_4152_));
 sky130_fd_sc_hd__buf_1 _8348_ (.A(_4152_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_2 _8349_ (.A0(\rf.registers[16][18] ),
    .A1(_3493_),
    .S(_4144_),
    .X(_4153_));
 sky130_fd_sc_hd__buf_1 _8350_ (.A(_4153_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_2 _8351_ (.A0(\rf.registers[16][19] ),
    .A1(_3495_),
    .S(_4144_),
    .X(_4154_));
 sky130_fd_sc_hd__buf_1 _8352_ (.A(_4154_),
    .X(_0649_));
 sky130_fd_sc_hd__buf_1 _8353_ (.A(_4132_),
    .X(_4155_));
 sky130_fd_sc_hd__mux2_2 _8354_ (.A0(\rf.registers[16][20] ),
    .A1(_3497_),
    .S(_4155_),
    .X(_4156_));
 sky130_fd_sc_hd__buf_1 _8355_ (.A(_4156_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_2 _8356_ (.A0(\rf.registers[16][21] ),
    .A1(_3500_),
    .S(_4155_),
    .X(_4157_));
 sky130_fd_sc_hd__buf_1 _8357_ (.A(_4157_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_2 _8358_ (.A0(\rf.registers[16][22] ),
    .A1(_3502_),
    .S(_4155_),
    .X(_4158_));
 sky130_fd_sc_hd__buf_1 _8359_ (.A(_4158_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_2 _8360_ (.A0(\rf.registers[16][23] ),
    .A1(_3504_),
    .S(_4155_),
    .X(_4159_));
 sky130_fd_sc_hd__buf_1 _8361_ (.A(_4159_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_2 _8362_ (.A0(\rf.registers[16][24] ),
    .A1(_3506_),
    .S(_4155_),
    .X(_4160_));
 sky130_fd_sc_hd__buf_1 _8363_ (.A(_4160_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_2 _8364_ (.A0(\rf.registers[16][25] ),
    .A1(_3508_),
    .S(_4155_),
    .X(_4161_));
 sky130_fd_sc_hd__buf_1 _8365_ (.A(_4161_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_2 _8366_ (.A0(\rf.registers[16][26] ),
    .A1(_3442_),
    .S(_4155_),
    .X(_4162_));
 sky130_fd_sc_hd__buf_1 _8367_ (.A(_4162_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_2 _8368_ (.A0(\rf.registers[16][27] ),
    .A1(_3444_),
    .S(_4155_),
    .X(_4163_));
 sky130_fd_sc_hd__buf_1 _8369_ (.A(_4163_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_2 _8370_ (.A0(\rf.registers[16][28] ),
    .A1(_3446_),
    .S(_4155_),
    .X(_4164_));
 sky130_fd_sc_hd__buf_1 _8371_ (.A(_4164_),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_2 _8372_ (.A0(\rf.registers[16][29] ),
    .A1(_3448_),
    .S(_4155_),
    .X(_4165_));
 sky130_fd_sc_hd__buf_1 _8373_ (.A(_4165_),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_2 _8374_ (.A0(\rf.registers[16][30] ),
    .A1(_3450_),
    .S(_4132_),
    .X(_4166_));
 sky130_fd_sc_hd__buf_1 _8375_ (.A(_4166_),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_2 _8376_ (.A0(\rf.registers[16][31] ),
    .A1(_3452_),
    .S(_4132_),
    .X(_4167_));
 sky130_fd_sc_hd__buf_1 _8377_ (.A(_4167_),
    .X(_0661_));
 sky130_fd_sc_hd__nor2b_2 _8378_ (.A(_3155_),
    .B_N(_3192_),
    .Y(_4168_));
 sky130_fd_sc_hd__buf_1 _8379_ (.A(_4168_),
    .X(_4169_));
 sky130_fd_sc_hd__mux2_2 _8380_ (.A0(\rf.registers[12][0] ),
    .A1(_3454_),
    .S(_4169_),
    .X(_4170_));
 sky130_fd_sc_hd__buf_1 _8381_ (.A(_4170_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_2 _8382_ (.A0(\rf.registers[12][1] ),
    .A1(_3458_),
    .S(_4169_),
    .X(_4171_));
 sky130_fd_sc_hd__buf_1 _8383_ (.A(_4171_),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_2 _8384_ (.A0(\rf.registers[12][2] ),
    .A1(_3460_),
    .S(_4169_),
    .X(_4172_));
 sky130_fd_sc_hd__buf_1 _8385_ (.A(_4172_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_2 _8386_ (.A0(\rf.registers[12][3] ),
    .A1(_3462_),
    .S(_4169_),
    .X(_4173_));
 sky130_fd_sc_hd__buf_1 _8387_ (.A(_4173_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_2 _8388_ (.A0(\rf.registers[12][4] ),
    .A1(_3464_),
    .S(_4169_),
    .X(_4174_));
 sky130_fd_sc_hd__buf_1 _8389_ (.A(_4174_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_2 _8390_ (.A0(\rf.registers[12][5] ),
    .A1(_3466_),
    .S(_4169_),
    .X(_4175_));
 sky130_fd_sc_hd__buf_1 _8391_ (.A(_4175_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_2 _8392_ (.A0(\rf.registers[12][6] ),
    .A1(_3468_),
    .S(_4169_),
    .X(_4176_));
 sky130_fd_sc_hd__buf_1 _8393_ (.A(_4176_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_2 _8394_ (.A0(\rf.registers[12][7] ),
    .A1(_3470_),
    .S(_4169_),
    .X(_4177_));
 sky130_fd_sc_hd__buf_1 _8395_ (.A(_4177_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_2 _8396_ (.A0(\rf.registers[12][8] ),
    .A1(_3472_),
    .S(_4169_),
    .X(_4178_));
 sky130_fd_sc_hd__buf_1 _8397_ (.A(_4178_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_2 _8398_ (.A0(\rf.registers[12][9] ),
    .A1(_3474_),
    .S(_4169_),
    .X(_4179_));
 sky130_fd_sc_hd__buf_1 _8399_ (.A(_4179_),
    .X(_0671_));
 sky130_fd_sc_hd__buf_1 _8400_ (.A(_4168_),
    .X(_4180_));
 sky130_fd_sc_hd__mux2_2 _8401_ (.A0(\rf.registers[12][10] ),
    .A1(_3476_),
    .S(_4180_),
    .X(_4181_));
 sky130_fd_sc_hd__buf_1 _8402_ (.A(_4181_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_2 _8403_ (.A0(\rf.registers[12][11] ),
    .A1(_3479_),
    .S(_4180_),
    .X(_4182_));
 sky130_fd_sc_hd__buf_1 _8404_ (.A(_4182_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_2 _8405_ (.A0(\rf.registers[12][12] ),
    .A1(_3481_),
    .S(_4180_),
    .X(_4183_));
 sky130_fd_sc_hd__buf_1 _8406_ (.A(_4183_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_2 _8407_ (.A0(\rf.registers[12][13] ),
    .A1(_3483_),
    .S(_4180_),
    .X(_4184_));
 sky130_fd_sc_hd__buf_1 _8408_ (.A(_4184_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_2 _8409_ (.A0(\rf.registers[12][14] ),
    .A1(_3485_),
    .S(_4180_),
    .X(_4185_));
 sky130_fd_sc_hd__buf_1 _8410_ (.A(_4185_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_2 _8411_ (.A0(\rf.registers[12][15] ),
    .A1(_3487_),
    .S(_4180_),
    .X(_4186_));
 sky130_fd_sc_hd__buf_1 _8412_ (.A(_4186_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_2 _8413_ (.A0(\rf.registers[12][16] ),
    .A1(_3489_),
    .S(_4180_),
    .X(_4187_));
 sky130_fd_sc_hd__buf_1 _8414_ (.A(_4187_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_2 _8415_ (.A0(\rf.registers[12][17] ),
    .A1(_3491_),
    .S(_4180_),
    .X(_4188_));
 sky130_fd_sc_hd__buf_1 _8416_ (.A(_4188_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_2 _8417_ (.A0(\rf.registers[12][18] ),
    .A1(_3493_),
    .S(_4180_),
    .X(_4189_));
 sky130_fd_sc_hd__buf_1 _8418_ (.A(_4189_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_2 _8419_ (.A0(\rf.registers[12][19] ),
    .A1(_3495_),
    .S(_4180_),
    .X(_4190_));
 sky130_fd_sc_hd__buf_1 _8420_ (.A(_4190_),
    .X(_0681_));
 sky130_fd_sc_hd__buf_1 _8421_ (.A(_4168_),
    .X(_4191_));
 sky130_fd_sc_hd__mux2_2 _8422_ (.A0(\rf.registers[12][20] ),
    .A1(_3497_),
    .S(_4191_),
    .X(_4192_));
 sky130_fd_sc_hd__buf_1 _8423_ (.A(_4192_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_2 _8424_ (.A0(\rf.registers[12][21] ),
    .A1(_3500_),
    .S(_4191_),
    .X(_4193_));
 sky130_fd_sc_hd__buf_1 _8425_ (.A(_4193_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_2 _8426_ (.A0(\rf.registers[12][22] ),
    .A1(_3502_),
    .S(_4191_),
    .X(_4194_));
 sky130_fd_sc_hd__buf_1 _8427_ (.A(_4194_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_2 _8428_ (.A0(\rf.registers[12][23] ),
    .A1(_3504_),
    .S(_4191_),
    .X(_4195_));
 sky130_fd_sc_hd__buf_1 _8429_ (.A(_4195_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_2 _8430_ (.A0(\rf.registers[12][24] ),
    .A1(_3506_),
    .S(_4191_),
    .X(_4196_));
 sky130_fd_sc_hd__buf_1 _8431_ (.A(_4196_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_2 _8432_ (.A0(\rf.registers[12][25] ),
    .A1(_3508_),
    .S(_4191_),
    .X(_4197_));
 sky130_fd_sc_hd__buf_1 _8433_ (.A(_4197_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_2 _8434_ (.A0(\rf.registers[12][26] ),
    .A1(WD3[26]),
    .S(_4191_),
    .X(_4198_));
 sky130_fd_sc_hd__buf_1 _8435_ (.A(_4198_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_2 _8436_ (.A0(\rf.registers[12][27] ),
    .A1(WD3[27]),
    .S(_4191_),
    .X(_4199_));
 sky130_fd_sc_hd__buf_1 _8437_ (.A(_4199_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_2 _8438_ (.A0(\rf.registers[12][28] ),
    .A1(WD3[28]),
    .S(_4191_),
    .X(_4200_));
 sky130_fd_sc_hd__buf_1 _8439_ (.A(_4200_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_2 _8440_ (.A0(\rf.registers[12][29] ),
    .A1(WD3[29]),
    .S(_4191_),
    .X(_4201_));
 sky130_fd_sc_hd__buf_1 _8441_ (.A(_4201_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_2 _8442_ (.A0(\rf.registers[12][30] ),
    .A1(WD3[30]),
    .S(_4168_),
    .X(_4202_));
 sky130_fd_sc_hd__buf_1 _8443_ (.A(_4202_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_2 _8444_ (.A0(\rf.registers[12][31] ),
    .A1(WD3[31]),
    .S(_4168_),
    .X(_4203_));
 sky130_fd_sc_hd__buf_1 _8445_ (.A(_4203_),
    .X(_0693_));
 sky130_fd_sc_hd__nor2_2 _8446_ (.A(_3003_),
    .B(_3411_),
    .Y(_4204_));
 sky130_fd_sc_hd__buf_1 _8447_ (.A(_4204_),
    .X(_4205_));
 sky130_fd_sc_hd__mux2_2 _8448_ (.A0(\rf.registers[11][0] ),
    .A1(WD3[0]),
    .S(_4205_),
    .X(_4206_));
 sky130_fd_sc_hd__buf_1 _8449_ (.A(_4206_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_2 _8450_ (.A0(\rf.registers[11][1] ),
    .A1(WD3[1]),
    .S(_4205_),
    .X(_4207_));
 sky130_fd_sc_hd__buf_1 _8451_ (.A(_4207_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_2 _8452_ (.A0(\rf.registers[11][2] ),
    .A1(WD3[2]),
    .S(_4205_),
    .X(_4208_));
 sky130_fd_sc_hd__buf_1 _8453_ (.A(_4208_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_2 _8454_ (.A0(\rf.registers[11][3] ),
    .A1(WD3[3]),
    .S(_4205_),
    .X(_4209_));
 sky130_fd_sc_hd__buf_1 _8455_ (.A(_4209_),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_2 _8456_ (.A0(\rf.registers[11][4] ),
    .A1(WD3[4]),
    .S(_4205_),
    .X(_4210_));
 sky130_fd_sc_hd__buf_1 _8457_ (.A(_4210_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_2 _8458_ (.A0(\rf.registers[11][5] ),
    .A1(WD3[5]),
    .S(_4205_),
    .X(_4211_));
 sky130_fd_sc_hd__buf_1 _8459_ (.A(_4211_),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_2 _8460_ (.A0(\rf.registers[11][6] ),
    .A1(WD3[6]),
    .S(_4205_),
    .X(_4212_));
 sky130_fd_sc_hd__buf_1 _8461_ (.A(_4212_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_2 _8462_ (.A0(\rf.registers[11][7] ),
    .A1(WD3[7]),
    .S(_4205_),
    .X(_4213_));
 sky130_fd_sc_hd__buf_1 _8463_ (.A(_4213_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_2 _8464_ (.A0(\rf.registers[11][8] ),
    .A1(WD3[8]),
    .S(_4205_),
    .X(_4214_));
 sky130_fd_sc_hd__buf_1 _8465_ (.A(_4214_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_2 _8466_ (.A0(\rf.registers[11][9] ),
    .A1(WD3[9]),
    .S(_4205_),
    .X(_4215_));
 sky130_fd_sc_hd__buf_1 _8467_ (.A(_4215_),
    .X(_0703_));
 sky130_fd_sc_hd__buf_1 _8468_ (.A(_4204_),
    .X(_4216_));
 sky130_fd_sc_hd__mux2_2 _8469_ (.A0(\rf.registers[11][10] ),
    .A1(WD3[10]),
    .S(_4216_),
    .X(_4217_));
 sky130_fd_sc_hd__buf_1 _8470_ (.A(_4217_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_2 _8471_ (.A0(\rf.registers[11][11] ),
    .A1(WD3[11]),
    .S(_4216_),
    .X(_4218_));
 sky130_fd_sc_hd__buf_1 _8472_ (.A(_4218_),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_2 _8473_ (.A0(\rf.registers[11][12] ),
    .A1(WD3[12]),
    .S(_4216_),
    .X(_4219_));
 sky130_fd_sc_hd__buf_1 _8474_ (.A(_4219_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_2 _8475_ (.A0(\rf.registers[11][13] ),
    .A1(WD3[13]),
    .S(_4216_),
    .X(_4220_));
 sky130_fd_sc_hd__buf_1 _8476_ (.A(_4220_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_2 _8477_ (.A0(\rf.registers[11][14] ),
    .A1(WD3[14]),
    .S(_4216_),
    .X(_4221_));
 sky130_fd_sc_hd__buf_1 _8478_ (.A(_4221_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_2 _8479_ (.A0(\rf.registers[11][15] ),
    .A1(WD3[15]),
    .S(_4216_),
    .X(_4222_));
 sky130_fd_sc_hd__buf_1 _8480_ (.A(_4222_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_2 _8481_ (.A0(\rf.registers[11][16] ),
    .A1(WD3[16]),
    .S(_4216_),
    .X(_4223_));
 sky130_fd_sc_hd__buf_1 _8482_ (.A(_4223_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_2 _8483_ (.A0(\rf.registers[11][17] ),
    .A1(WD3[17]),
    .S(_4216_),
    .X(_4224_));
 sky130_fd_sc_hd__buf_1 _8484_ (.A(_4224_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_2 _8485_ (.A0(\rf.registers[11][18] ),
    .A1(WD3[18]),
    .S(_4216_),
    .X(_4225_));
 sky130_fd_sc_hd__buf_1 _8486_ (.A(_4225_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_2 _8487_ (.A0(\rf.registers[11][19] ),
    .A1(WD3[19]),
    .S(_4216_),
    .X(_4226_));
 sky130_fd_sc_hd__buf_1 _8488_ (.A(_4226_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_1 _8489_ (.A(_4204_),
    .X(_4227_));
 sky130_fd_sc_hd__mux2_2 _8490_ (.A0(\rf.registers[11][20] ),
    .A1(WD3[20]),
    .S(_4227_),
    .X(_4228_));
 sky130_fd_sc_hd__buf_1 _8491_ (.A(_4228_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_2 _8492_ (.A0(\rf.registers[11][21] ),
    .A1(WD3[21]),
    .S(_4227_),
    .X(_4229_));
 sky130_fd_sc_hd__buf_1 _8493_ (.A(_4229_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_2 _8494_ (.A0(\rf.registers[11][22] ),
    .A1(WD3[22]),
    .S(_4227_),
    .X(_4230_));
 sky130_fd_sc_hd__buf_1 _8495_ (.A(_4230_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_2 _8496_ (.A0(\rf.registers[11][23] ),
    .A1(WD3[23]),
    .S(_4227_),
    .X(_4231_));
 sky130_fd_sc_hd__buf_1 _8497_ (.A(_4231_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_2 _8498_ (.A0(\rf.registers[11][24] ),
    .A1(WD3[24]),
    .S(_4227_),
    .X(_4232_));
 sky130_fd_sc_hd__buf_1 _8499_ (.A(_4232_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_2 _8500_ (.A0(\rf.registers[11][25] ),
    .A1(WD3[25]),
    .S(_4227_),
    .X(_4233_));
 sky130_fd_sc_hd__buf_1 _8501_ (.A(_4233_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_2 _8502_ (.A0(\rf.registers[11][26] ),
    .A1(WD3[26]),
    .S(_4227_),
    .X(_4234_));
 sky130_fd_sc_hd__buf_1 _8503_ (.A(_4234_),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_2 _8504_ (.A0(\rf.registers[11][27] ),
    .A1(WD3[27]),
    .S(_4227_),
    .X(_4235_));
 sky130_fd_sc_hd__buf_1 _8505_ (.A(_4235_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_2 _8506_ (.A0(\rf.registers[11][28] ),
    .A1(WD3[28]),
    .S(_4227_),
    .X(_4236_));
 sky130_fd_sc_hd__buf_1 _8507_ (.A(_4236_),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_2 _8508_ (.A0(\rf.registers[11][29] ),
    .A1(WD3[29]),
    .S(_4227_),
    .X(_4237_));
 sky130_fd_sc_hd__buf_1 _8509_ (.A(_4237_),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_2 _8510_ (.A0(\rf.registers[11][30] ),
    .A1(WD3[30]),
    .S(_4204_),
    .X(_4238_));
 sky130_fd_sc_hd__buf_1 _8511_ (.A(_4238_),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_2 _8512_ (.A0(\rf.registers[11][31] ),
    .A1(WD3[31]),
    .S(_4204_),
    .X(_4239_));
 sky130_fd_sc_hd__buf_1 _8513_ (.A(_4239_),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_2 _8514_ (.A0(\rf.registers[10][0] ),
    .A1(WD3[0]),
    .S(_3007_),
    .X(_4240_));
 sky130_fd_sc_hd__buf_1 _8515_ (.A(_4240_),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_2 _8516_ (.A0(\rf.registers[10][1] ),
    .A1(WD3[1]),
    .S(_3007_),
    .X(_4241_));
 sky130_fd_sc_hd__buf_1 _8517_ (.A(_4241_),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_2 _8518_ (.A0(\rf.registers[10][2] ),
    .A1(WD3[2]),
    .S(_3007_),
    .X(_4242_));
 sky130_fd_sc_hd__buf_1 _8519_ (.A(_4242_),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_2 _8520_ (.A0(\rf.registers[10][3] ),
    .A1(WD3[3]),
    .S(_3007_),
    .X(_4243_));
 sky130_fd_sc_hd__buf_1 _8521_ (.A(_4243_),
    .X(_0729_));
 sky130_fd_sc_hd__buf_1 _8522_ (.A(_3006_),
    .X(_4244_));
 sky130_fd_sc_hd__mux2_2 _8523_ (.A0(\rf.registers[10][4] ),
    .A1(WD3[4]),
    .S(_4244_),
    .X(_4245_));
 sky130_fd_sc_hd__buf_1 _8524_ (.A(_4245_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_2 _8525_ (.A0(\rf.registers[10][5] ),
    .A1(WD3[5]),
    .S(_4244_),
    .X(_4246_));
 sky130_fd_sc_hd__buf_1 _8526_ (.A(_4246_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_2 _8527_ (.A0(\rf.registers[10][6] ),
    .A1(WD3[6]),
    .S(_4244_),
    .X(_4247_));
 sky130_fd_sc_hd__buf_1 _8528_ (.A(_4247_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_2 _8529_ (.A0(\rf.registers[10][7] ),
    .A1(WD3[7]),
    .S(_4244_),
    .X(_4248_));
 sky130_fd_sc_hd__buf_1 _8530_ (.A(_4248_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_2 _8531_ (.A0(\rf.registers[10][8] ),
    .A1(WD3[8]),
    .S(_4244_),
    .X(_4249_));
 sky130_fd_sc_hd__buf_1 _8532_ (.A(_4249_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_2 _8533_ (.A0(\rf.registers[10][9] ),
    .A1(WD3[9]),
    .S(_4244_),
    .X(_4250_));
 sky130_fd_sc_hd__buf_1 _8534_ (.A(_4250_),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_2 _8535_ (.A0(\rf.registers[10][10] ),
    .A1(WD3[10]),
    .S(_4244_),
    .X(_4251_));
 sky130_fd_sc_hd__buf_1 _8536_ (.A(_4251_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_2 _8537_ (.A0(\rf.registers[10][11] ),
    .A1(WD3[11]),
    .S(_4244_),
    .X(_4252_));
 sky130_fd_sc_hd__buf_1 _8538_ (.A(_4252_),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_2 _8539_ (.A0(\rf.registers[10][12] ),
    .A1(WD3[12]),
    .S(_4244_),
    .X(_4253_));
 sky130_fd_sc_hd__buf_1 _8540_ (.A(_4253_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_2 _8541_ (.A0(\rf.registers[10][13] ),
    .A1(WD3[13]),
    .S(_4244_),
    .X(_4254_));
 sky130_fd_sc_hd__buf_1 _8542_ (.A(_4254_),
    .X(_0739_));
 sky130_fd_sc_hd__buf_1 _8543_ (.A(_3006_),
    .X(_4255_));
 sky130_fd_sc_hd__mux2_2 _8544_ (.A0(\rf.registers[10][14] ),
    .A1(WD3[14]),
    .S(_4255_),
    .X(_4256_));
 sky130_fd_sc_hd__buf_1 _8545_ (.A(_4256_),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_2 _8546_ (.A0(\rf.registers[10][15] ),
    .A1(WD3[15]),
    .S(_4255_),
    .X(_4257_));
 sky130_fd_sc_hd__buf_1 _8547_ (.A(_4257_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_2 _8548_ (.A0(\rf.registers[10][16] ),
    .A1(WD3[16]),
    .S(_4255_),
    .X(_4258_));
 sky130_fd_sc_hd__buf_1 _8549_ (.A(_4258_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_2 _8550_ (.A0(\rf.registers[10][17] ),
    .A1(WD3[17]),
    .S(_4255_),
    .X(_4259_));
 sky130_fd_sc_hd__buf_1 _8551_ (.A(_4259_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_2 _8552_ (.A0(\rf.registers[10][18] ),
    .A1(WD3[18]),
    .S(_4255_),
    .X(_4260_));
 sky130_fd_sc_hd__buf_1 _8553_ (.A(_4260_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_2 _8554_ (.A0(\rf.registers[10][19] ),
    .A1(WD3[19]),
    .S(_4255_),
    .X(_4261_));
 sky130_fd_sc_hd__buf_1 _8555_ (.A(_4261_),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_2 _8556_ (.A0(\rf.registers[10][20] ),
    .A1(WD3[20]),
    .S(_4255_),
    .X(_4262_));
 sky130_fd_sc_hd__buf_1 _8557_ (.A(_4262_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_2 _8558_ (.A0(\rf.registers[10][21] ),
    .A1(WD3[21]),
    .S(_4255_),
    .X(_4263_));
 sky130_fd_sc_hd__buf_1 _8559_ (.A(_4263_),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_2 _8560_ (.A0(\rf.registers[10][22] ),
    .A1(WD3[22]),
    .S(_4255_),
    .X(_4264_));
 sky130_fd_sc_hd__buf_1 _8561_ (.A(_4264_),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_2 _8562_ (.A0(\rf.registers[10][23] ),
    .A1(WD3[23]),
    .S(_4255_),
    .X(_4265_));
 sky130_fd_sc_hd__buf_1 _8563_ (.A(_4265_),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_2 _8564_ (.A0(\rf.registers[10][24] ),
    .A1(WD3[24]),
    .S(_3006_),
    .X(_4266_));
 sky130_fd_sc_hd__buf_1 _8565_ (.A(_4266_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_2 _8566_ (.A0(\rf.registers[10][25] ),
    .A1(WD3[25]),
    .S(_3006_),
    .X(_4267_));
 sky130_fd_sc_hd__buf_1 _8567_ (.A(_4267_),
    .X(_0751_));
 sky130_fd_sc_hd__dfxtp_2 _8568_ (.CLK(clk),
    .D(_0752_),
    .Q(\rf.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8569_ (.CLK(clk),
    .D(_0753_),
    .Q(\rf.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8570_ (.CLK(clk),
    .D(_0754_),
    .Q(\rf.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8571_ (.CLK(clk),
    .D(_0755_),
    .Q(\rf.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8572_ (.CLK(clk),
    .D(_0756_),
    .Q(\rf.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8573_ (.CLK(clk),
    .D(_0757_),
    .Q(\rf.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8574_ (.CLK(clk),
    .D(_0758_),
    .Q(\rf.registers[22][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8575_ (.CLK(clk),
    .D(_0759_),
    .Q(\rf.registers[22][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8576_ (.CLK(clk),
    .D(_0760_),
    .Q(\rf.registers[22][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8577_ (.CLK(clk),
    .D(_0761_),
    .Q(\rf.registers[22][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8578_ (.CLK(clk),
    .D(_0762_),
    .Q(\rf.registers[22][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8579_ (.CLK(clk),
    .D(_0763_),
    .Q(\rf.registers[22][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8580_ (.CLK(clk),
    .D(_0764_),
    .Q(\rf.registers[22][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8581_ (.CLK(clk),
    .D(_0765_),
    .Q(\rf.registers[22][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8582_ (.CLK(clk),
    .D(_0766_),
    .Q(\rf.registers[22][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8583_ (.CLK(clk),
    .D(_0767_),
    .Q(\rf.registers[22][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8584_ (.CLK(clk),
    .D(_0768_),
    .Q(\rf.registers[22][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8585_ (.CLK(clk),
    .D(_0769_),
    .Q(\rf.registers[22][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8586_ (.CLK(clk),
    .D(_0770_),
    .Q(\rf.registers[22][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8587_ (.CLK(clk),
    .D(_0771_),
    .Q(\rf.registers[22][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8588_ (.CLK(clk),
    .D(_0772_),
    .Q(\rf.registers[22][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8589_ (.CLK(clk),
    .D(_0773_),
    .Q(\rf.registers[22][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8590_ (.CLK(clk),
    .D(_0774_),
    .Q(\rf.registers[22][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8591_ (.CLK(clk),
    .D(_0775_),
    .Q(\rf.registers[22][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8592_ (.CLK(clk),
    .D(_0776_),
    .Q(\rf.registers[22][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8593_ (.CLK(clk),
    .D(_0777_),
    .Q(\rf.registers[22][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8594_ (.CLK(clk),
    .D(_0778_),
    .Q(\rf.registers[22][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8595_ (.CLK(clk),
    .D(_0779_),
    .Q(\rf.registers[22][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8596_ (.CLK(clk),
    .D(_0780_),
    .Q(\rf.registers[22][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8597_ (.CLK(clk),
    .D(_0781_),
    .Q(\rf.registers[22][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8598_ (.CLK(clk),
    .D(_0782_),
    .Q(\rf.registers[22][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8599_ (.CLK(clk),
    .D(_0783_),
    .Q(\rf.registers[22][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8600_ (.CLK(clk),
    .D(_0784_),
    .Q(\rf.registers[22][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8601_ (.CLK(clk),
    .D(_0785_),
    .Q(\rf.registers[22][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8602_ (.CLK(clk),
    .D(_0786_),
    .Q(\rf.registers[22][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8603_ (.CLK(clk),
    .D(_0787_),
    .Q(\rf.registers[22][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8604_ (.CLK(clk),
    .D(_0788_),
    .Q(\rf.registers[22][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8605_ (.CLK(clk),
    .D(_0789_),
    .Q(\rf.registers[22][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8606_ (.CLK(clk),
    .D(_0790_),
    .Q(\rf.registers[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8607_ (.CLK(clk),
    .D(_0791_),
    .Q(\rf.registers[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8608_ (.CLK(clk),
    .D(_0792_),
    .Q(\rf.registers[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8609_ (.CLK(clk),
    .D(_0793_),
    .Q(\rf.registers[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8610_ (.CLK(clk),
    .D(_0794_),
    .Q(\rf.registers[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8611_ (.CLK(clk),
    .D(_0795_),
    .Q(\rf.registers[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8612_ (.CLK(clk),
    .D(_0796_),
    .Q(\rf.registers[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8613_ (.CLK(clk),
    .D(_0797_),
    .Q(\rf.registers[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8614_ (.CLK(clk),
    .D(_0798_),
    .Q(\rf.registers[17][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8615_ (.CLK(clk),
    .D(_0799_),
    .Q(\rf.registers[17][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8616_ (.CLK(clk),
    .D(_0800_),
    .Q(\rf.registers[17][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8617_ (.CLK(clk),
    .D(_0801_),
    .Q(\rf.registers[17][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8618_ (.CLK(clk),
    .D(_0802_),
    .Q(\rf.registers[17][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8619_ (.CLK(clk),
    .D(_0803_),
    .Q(\rf.registers[17][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8620_ (.CLK(clk),
    .D(_0804_),
    .Q(\rf.registers[17][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8621_ (.CLK(clk),
    .D(_0805_),
    .Q(\rf.registers[17][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8622_ (.CLK(clk),
    .D(_0806_),
    .Q(\rf.registers[17][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8623_ (.CLK(clk),
    .D(_0807_),
    .Q(\rf.registers[17][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8624_ (.CLK(clk),
    .D(_0808_),
    .Q(\rf.registers[17][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8625_ (.CLK(clk),
    .D(_0809_),
    .Q(\rf.registers[17][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8626_ (.CLK(clk),
    .D(_0810_),
    .Q(\rf.registers[17][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8627_ (.CLK(clk),
    .D(_0811_),
    .Q(\rf.registers[17][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8628_ (.CLK(clk),
    .D(_0812_),
    .Q(\rf.registers[17][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8629_ (.CLK(clk),
    .D(_0813_),
    .Q(\rf.registers[17][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8630_ (.CLK(clk),
    .D(_0814_),
    .Q(\rf.registers[17][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8631_ (.CLK(clk),
    .D(_0815_),
    .Q(\rf.registers[17][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8632_ (.CLK(clk),
    .D(_0816_),
    .Q(\rf.registers[17][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8633_ (.CLK(clk),
    .D(_0817_),
    .Q(\rf.registers[17][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8634_ (.CLK(clk),
    .D(_0818_),
    .Q(\rf.registers[17][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8635_ (.CLK(clk),
    .D(_0819_),
    .Q(\rf.registers[17][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8636_ (.CLK(clk),
    .D(_0820_),
    .Q(\rf.registers[17][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8637_ (.CLK(clk),
    .D(_0821_),
    .Q(\rf.registers[17][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8638_ (.CLK(clk),
    .D(_0822_),
    .Q(\rf.registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8639_ (.CLK(clk),
    .D(_0823_),
    .Q(\rf.registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8640_ (.CLK(clk),
    .D(_0824_),
    .Q(\rf.registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8641_ (.CLK(clk),
    .D(_0825_),
    .Q(\rf.registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8642_ (.CLK(clk),
    .D(_0826_),
    .Q(\rf.registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8643_ (.CLK(clk),
    .D(_0827_),
    .Q(\rf.registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8644_ (.CLK(clk),
    .D(_0828_),
    .Q(\rf.registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8645_ (.CLK(clk),
    .D(_0829_),
    .Q(\rf.registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8646_ (.CLK(clk),
    .D(_0830_),
    .Q(\rf.registers[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8647_ (.CLK(clk),
    .D(_0831_),
    .Q(\rf.registers[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8648_ (.CLK(clk),
    .D(_0832_),
    .Q(\rf.registers[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8649_ (.CLK(clk),
    .D(_0833_),
    .Q(\rf.registers[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8650_ (.CLK(clk),
    .D(_0834_),
    .Q(\rf.registers[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8651_ (.CLK(clk),
    .D(_0835_),
    .Q(\rf.registers[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8652_ (.CLK(clk),
    .D(_0836_),
    .Q(\rf.registers[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8653_ (.CLK(clk),
    .D(_0837_),
    .Q(\rf.registers[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8654_ (.CLK(clk),
    .D(_0838_),
    .Q(\rf.registers[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8655_ (.CLK(clk),
    .D(_0839_),
    .Q(\rf.registers[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8656_ (.CLK(clk),
    .D(_0840_),
    .Q(\rf.registers[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8657_ (.CLK(clk),
    .D(_0841_),
    .Q(\rf.registers[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8658_ (.CLK(clk),
    .D(_0842_),
    .Q(\rf.registers[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8659_ (.CLK(clk),
    .D(_0843_),
    .Q(\rf.registers[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8660_ (.CLK(clk),
    .D(_0844_),
    .Q(\rf.registers[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8661_ (.CLK(clk),
    .D(_0845_),
    .Q(\rf.registers[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8662_ (.CLK(clk),
    .D(_0846_),
    .Q(\rf.registers[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8663_ (.CLK(clk),
    .D(_0847_),
    .Q(\rf.registers[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8664_ (.CLK(clk),
    .D(_0848_),
    .Q(\rf.registers[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8665_ (.CLK(clk),
    .D(_0849_),
    .Q(\rf.registers[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8666_ (.CLK(clk),
    .D(_0850_),
    .Q(\rf.registers[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8667_ (.CLK(clk),
    .D(_0851_),
    .Q(\rf.registers[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8668_ (.CLK(clk),
    .D(_0852_),
    .Q(\rf.registers[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8669_ (.CLK(clk),
    .D(_0853_),
    .Q(\rf.registers[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8670_ (.CLK(clk),
    .D(_0854_),
    .Q(\rf.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8671_ (.CLK(clk),
    .D(_0855_),
    .Q(\rf.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8672_ (.CLK(clk),
    .D(_0856_),
    .Q(\rf.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8673_ (.CLK(clk),
    .D(_0857_),
    .Q(\rf.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8674_ (.CLK(clk),
    .D(_0858_),
    .Q(\rf.registers[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8675_ (.CLK(clk),
    .D(_0859_),
    .Q(\rf.registers[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8676_ (.CLK(clk),
    .D(_0860_),
    .Q(\rf.registers[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8677_ (.CLK(clk),
    .D(_0861_),
    .Q(\rf.registers[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8678_ (.CLK(clk),
    .D(_0862_),
    .Q(\rf.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8679_ (.CLK(clk),
    .D(_0863_),
    .Q(\rf.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8680_ (.CLK(clk),
    .D(_0864_),
    .Q(\rf.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8681_ (.CLK(clk),
    .D(_0865_),
    .Q(\rf.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8682_ (.CLK(clk),
    .D(_0866_),
    .Q(\rf.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8683_ (.CLK(clk),
    .D(_0867_),
    .Q(\rf.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8684_ (.CLK(clk),
    .D(_0868_),
    .Q(\rf.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8685_ (.CLK(clk),
    .D(_0869_),
    .Q(\rf.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8686_ (.CLK(clk),
    .D(_0870_),
    .Q(\rf.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8687_ (.CLK(clk),
    .D(_0871_),
    .Q(\rf.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8688_ (.CLK(clk),
    .D(_0872_),
    .Q(\rf.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8689_ (.CLK(clk),
    .D(_0873_),
    .Q(\rf.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8690_ (.CLK(clk),
    .D(_0874_),
    .Q(\rf.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8691_ (.CLK(clk),
    .D(_0875_),
    .Q(\rf.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8692_ (.CLK(clk),
    .D(_0876_),
    .Q(\rf.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8693_ (.CLK(clk),
    .D(_0877_),
    .Q(\rf.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8694_ (.CLK(clk),
    .D(_0878_),
    .Q(\rf.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8695_ (.CLK(clk),
    .D(_0879_),
    .Q(\rf.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8696_ (.CLK(clk),
    .D(_0880_),
    .Q(\rf.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8697_ (.CLK(clk),
    .D(_0881_),
    .Q(\rf.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8698_ (.CLK(clk),
    .D(_0882_),
    .Q(\rf.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8699_ (.CLK(clk),
    .D(_0883_),
    .Q(\rf.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8700_ (.CLK(clk),
    .D(_0884_),
    .Q(\rf.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8701_ (.CLK(clk),
    .D(_0885_),
    .Q(\rf.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8702_ (.CLK(clk),
    .D(_0886_),
    .Q(\rf.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8703_ (.CLK(clk),
    .D(_0887_),
    .Q(\rf.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8704_ (.CLK(clk),
    .D(_0888_),
    .Q(\rf.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8705_ (.CLK(clk),
    .D(_0889_),
    .Q(\rf.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8706_ (.CLK(clk),
    .D(_0890_),
    .Q(\rf.registers[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8707_ (.CLK(clk),
    .D(_0891_),
    .Q(\rf.registers[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8708_ (.CLK(clk),
    .D(_0892_),
    .Q(\rf.registers[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8709_ (.CLK(clk),
    .D(_0893_),
    .Q(\rf.registers[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8710_ (.CLK(clk),
    .D(_0894_),
    .Q(\rf.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8711_ (.CLK(clk),
    .D(_0895_),
    .Q(\rf.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8712_ (.CLK(clk),
    .D(_0896_),
    .Q(\rf.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8713_ (.CLK(clk),
    .D(_0897_),
    .Q(\rf.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8714_ (.CLK(clk),
    .D(_0898_),
    .Q(\rf.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8715_ (.CLK(clk),
    .D(_0899_),
    .Q(\rf.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8716_ (.CLK(clk),
    .D(_0900_),
    .Q(\rf.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8717_ (.CLK(clk),
    .D(_0901_),
    .Q(\rf.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8718_ (.CLK(clk),
    .D(_0902_),
    .Q(\rf.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8719_ (.CLK(clk),
    .D(_0903_),
    .Q(\rf.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8720_ (.CLK(clk),
    .D(_0904_),
    .Q(\rf.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8721_ (.CLK(clk),
    .D(_0905_),
    .Q(\rf.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8722_ (.CLK(clk),
    .D(_0906_),
    .Q(\rf.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8723_ (.CLK(clk),
    .D(_0907_),
    .Q(\rf.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8724_ (.CLK(clk),
    .D(_0908_),
    .Q(\rf.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8725_ (.CLK(clk),
    .D(_0909_),
    .Q(\rf.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8726_ (.CLK(clk),
    .D(_0910_),
    .Q(\rf.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8727_ (.CLK(clk),
    .D(_0911_),
    .Q(\rf.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8728_ (.CLK(clk),
    .D(_0912_),
    .Q(\rf.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8729_ (.CLK(clk),
    .D(_0913_),
    .Q(\rf.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8730_ (.CLK(clk),
    .D(_0914_),
    .Q(\rf.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8731_ (.CLK(clk),
    .D(_0915_),
    .Q(\rf.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8732_ (.CLK(clk),
    .D(_0916_),
    .Q(\rf.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8733_ (.CLK(clk),
    .D(_0917_),
    .Q(\rf.registers[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8734_ (.CLK(clk),
    .D(_0918_),
    .Q(\rf.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8735_ (.CLK(clk),
    .D(_0919_),
    .Q(\rf.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8736_ (.CLK(clk),
    .D(_0920_),
    .Q(\rf.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8737_ (.CLK(clk),
    .D(_0921_),
    .Q(\rf.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8738_ (.CLK(clk),
    .D(_0922_),
    .Q(\rf.registers[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8739_ (.CLK(clk),
    .D(_0923_),
    .Q(\rf.registers[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8740_ (.CLK(clk),
    .D(_0924_),
    .Q(\rf.registers[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8741_ (.CLK(clk),
    .D(_0925_),
    .Q(\rf.registers[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8742_ (.CLK(clk),
    .D(_0926_),
    .Q(\rf.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8743_ (.CLK(clk),
    .D(_0927_),
    .Q(\rf.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8744_ (.CLK(clk),
    .D(_0928_),
    .Q(\rf.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8745_ (.CLK(clk),
    .D(_0929_),
    .Q(\rf.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8746_ (.CLK(clk),
    .D(_0930_),
    .Q(\rf.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8747_ (.CLK(clk),
    .D(_0931_),
    .Q(\rf.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8748_ (.CLK(clk),
    .D(_0932_),
    .Q(\rf.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8749_ (.CLK(clk),
    .D(_0933_),
    .Q(\rf.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8750_ (.CLK(clk),
    .D(_0934_),
    .Q(\rf.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8751_ (.CLK(clk),
    .D(_0935_),
    .Q(\rf.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8752_ (.CLK(clk),
    .D(_0936_),
    .Q(\rf.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8753_ (.CLK(clk),
    .D(_0937_),
    .Q(\rf.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8754_ (.CLK(clk),
    .D(_0938_),
    .Q(\rf.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8755_ (.CLK(clk),
    .D(_0939_),
    .Q(\rf.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8756_ (.CLK(clk),
    .D(_0940_),
    .Q(\rf.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8757_ (.CLK(clk),
    .D(_0941_),
    .Q(\rf.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8758_ (.CLK(clk),
    .D(_0942_),
    .Q(\rf.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8759_ (.CLK(clk),
    .D(_0943_),
    .Q(\rf.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8760_ (.CLK(clk),
    .D(_0944_),
    .Q(\rf.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8761_ (.CLK(clk),
    .D(_0945_),
    .Q(\rf.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8762_ (.CLK(clk),
    .D(_0946_),
    .Q(\rf.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8763_ (.CLK(clk),
    .D(_0947_),
    .Q(\rf.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8764_ (.CLK(clk),
    .D(_0948_),
    .Q(\rf.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8765_ (.CLK(clk),
    .D(_0949_),
    .Q(\rf.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8766_ (.CLK(clk),
    .D(_0950_),
    .Q(\rf.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8767_ (.CLK(clk),
    .D(_0951_),
    .Q(\rf.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8768_ (.CLK(clk),
    .D(_0952_),
    .Q(\rf.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8769_ (.CLK(clk),
    .D(_0953_),
    .Q(\rf.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8770_ (.CLK(clk),
    .D(_0954_),
    .Q(\rf.registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8771_ (.CLK(clk),
    .D(_0955_),
    .Q(\rf.registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8772_ (.CLK(clk),
    .D(_0956_),
    .Q(\rf.registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8773_ (.CLK(clk),
    .D(_0957_),
    .Q(\rf.registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8774_ (.CLK(clk),
    .D(_0958_),
    .Q(\rf.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8775_ (.CLK(clk),
    .D(_0959_),
    .Q(\rf.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8776_ (.CLK(clk),
    .D(_0960_),
    .Q(\rf.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8777_ (.CLK(clk),
    .D(_0961_),
    .Q(\rf.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8778_ (.CLK(clk),
    .D(_0962_),
    .Q(\rf.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8779_ (.CLK(clk),
    .D(_0963_),
    .Q(\rf.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8780_ (.CLK(clk),
    .D(_0964_),
    .Q(\rf.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8781_ (.CLK(clk),
    .D(_0965_),
    .Q(\rf.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8782_ (.CLK(clk),
    .D(_0966_),
    .Q(\rf.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8783_ (.CLK(clk),
    .D(_0967_),
    .Q(\rf.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8784_ (.CLK(clk),
    .D(_0968_),
    .Q(\rf.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8785_ (.CLK(clk),
    .D(_0969_),
    .Q(\rf.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8786_ (.CLK(clk),
    .D(_0970_),
    .Q(\rf.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8787_ (.CLK(clk),
    .D(_0971_),
    .Q(\rf.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8788_ (.CLK(clk),
    .D(_0972_),
    .Q(\rf.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8789_ (.CLK(clk),
    .D(_0973_),
    .Q(\rf.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8790_ (.CLK(clk),
    .D(_0974_),
    .Q(\rf.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8791_ (.CLK(clk),
    .D(_0975_),
    .Q(\rf.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8792_ (.CLK(clk),
    .D(_0976_),
    .Q(\rf.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8793_ (.CLK(clk),
    .D(_0977_),
    .Q(\rf.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8794_ (.CLK(clk),
    .D(_0978_),
    .Q(\rf.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8795_ (.CLK(clk),
    .D(_0979_),
    .Q(\rf.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8796_ (.CLK(clk),
    .D(_0980_),
    .Q(\rf.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8797_ (.CLK(clk),
    .D(_0981_),
    .Q(\rf.registers[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8798_ (.CLK(clk),
    .D(_0982_),
    .Q(\rf.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8799_ (.CLK(clk),
    .D(_0983_),
    .Q(\rf.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8800_ (.CLK(clk),
    .D(_0984_),
    .Q(\rf.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8801_ (.CLK(clk),
    .D(_0985_),
    .Q(\rf.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8802_ (.CLK(clk),
    .D(_0986_),
    .Q(\rf.registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8803_ (.CLK(clk),
    .D(_0987_),
    .Q(\rf.registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8804_ (.CLK(clk),
    .D(_0988_),
    .Q(\rf.registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8805_ (.CLK(clk),
    .D(_0989_),
    .Q(\rf.registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8806_ (.CLK(clk),
    .D(_0990_),
    .Q(\rf.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8807_ (.CLK(clk),
    .D(_0991_),
    .Q(\rf.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8808_ (.CLK(clk),
    .D(_0992_),
    .Q(\rf.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8809_ (.CLK(clk),
    .D(_0993_),
    .Q(\rf.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8810_ (.CLK(clk),
    .D(_0994_),
    .Q(\rf.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8811_ (.CLK(clk),
    .D(_0995_),
    .Q(\rf.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8812_ (.CLK(clk),
    .D(_0996_),
    .Q(\rf.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8813_ (.CLK(clk),
    .D(_0997_),
    .Q(\rf.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8814_ (.CLK(clk),
    .D(_0998_),
    .Q(\rf.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8815_ (.CLK(clk),
    .D(_0999_),
    .Q(\rf.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8816_ (.CLK(clk),
    .D(_1000_),
    .Q(\rf.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8817_ (.CLK(clk),
    .D(_1001_),
    .Q(\rf.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8818_ (.CLK(clk),
    .D(_1002_),
    .Q(\rf.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8819_ (.CLK(clk),
    .D(_1003_),
    .Q(\rf.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8820_ (.CLK(clk),
    .D(_1004_),
    .Q(\rf.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8821_ (.CLK(clk),
    .D(_1005_),
    .Q(\rf.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8822_ (.CLK(clk),
    .D(_1006_),
    .Q(\rf.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8823_ (.CLK(clk),
    .D(_1007_),
    .Q(\rf.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8824_ (.CLK(clk),
    .D(_1008_),
    .Q(\rf.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8825_ (.CLK(clk),
    .D(_1009_),
    .Q(\rf.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8826_ (.CLK(clk),
    .D(_1010_),
    .Q(\rf.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8827_ (.CLK(clk),
    .D(_1011_),
    .Q(\rf.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8828_ (.CLK(clk),
    .D(_1012_),
    .Q(\rf.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8829_ (.CLK(clk),
    .D(_1013_),
    .Q(\rf.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8830_ (.CLK(clk),
    .D(_1014_),
    .Q(\rf.registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8831_ (.CLK(clk),
    .D(_1015_),
    .Q(\rf.registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8832_ (.CLK(clk),
    .D(_1016_),
    .Q(\rf.registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8833_ (.CLK(clk),
    .D(_1017_),
    .Q(\rf.registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8834_ (.CLK(clk),
    .D(_1018_),
    .Q(\rf.registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8835_ (.CLK(clk),
    .D(_1019_),
    .Q(\rf.registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8836_ (.CLK(clk),
    .D(_1020_),
    .Q(\rf.registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8837_ (.CLK(clk),
    .D(_1021_),
    .Q(\rf.registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8838_ (.CLK(clk),
    .D(_1022_),
    .Q(\rf.registers[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8839_ (.CLK(clk),
    .D(_1023_),
    .Q(\rf.registers[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8840_ (.CLK(clk),
    .D(_0000_),
    .Q(\rf.registers[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8841_ (.CLK(clk),
    .D(_0001_),
    .Q(\rf.registers[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8842_ (.CLK(clk),
    .D(_0002_),
    .Q(\rf.registers[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8843_ (.CLK(clk),
    .D(_0003_),
    .Q(\rf.registers[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8844_ (.CLK(clk),
    .D(_0004_),
    .Q(\rf.registers[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8845_ (.CLK(clk),
    .D(_0005_),
    .Q(\rf.registers[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8846_ (.CLK(clk),
    .D(_0006_),
    .Q(\rf.registers[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8847_ (.CLK(clk),
    .D(_0007_),
    .Q(\rf.registers[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8848_ (.CLK(clk),
    .D(_0008_),
    .Q(\rf.registers[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8849_ (.CLK(clk),
    .D(_0009_),
    .Q(\rf.registers[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8850_ (.CLK(clk),
    .D(_0010_),
    .Q(\rf.registers[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8851_ (.CLK(clk),
    .D(_0011_),
    .Q(\rf.registers[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8852_ (.CLK(clk),
    .D(_0012_),
    .Q(\rf.registers[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8853_ (.CLK(clk),
    .D(_0013_),
    .Q(\rf.registers[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8854_ (.CLK(clk),
    .D(_0014_),
    .Q(\rf.registers[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8855_ (.CLK(clk),
    .D(_0015_),
    .Q(\rf.registers[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8856_ (.CLK(clk),
    .D(_0016_),
    .Q(\rf.registers[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8857_ (.CLK(clk),
    .D(_0017_),
    .Q(\rf.registers[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8858_ (.CLK(clk),
    .D(_0018_),
    .Q(\rf.registers[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8859_ (.CLK(clk),
    .D(_0019_),
    .Q(\rf.registers[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8860_ (.CLK(clk),
    .D(_0020_),
    .Q(\rf.registers[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8861_ (.CLK(clk),
    .D(_0021_),
    .Q(\rf.registers[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8862_ (.CLK(clk),
    .D(_0022_),
    .Q(\rf.registers[19][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8863_ (.CLK(clk),
    .D(_0023_),
    .Q(\rf.registers[19][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8864_ (.CLK(clk),
    .D(_0024_),
    .Q(\rf.registers[19][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8865_ (.CLK(clk),
    .D(_0025_),
    .Q(\rf.registers[19][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8866_ (.CLK(clk),
    .D(_0026_),
    .Q(\rf.registers[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8867_ (.CLK(clk),
    .D(_0027_),
    .Q(\rf.registers[19][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8868_ (.CLK(clk),
    .D(_0028_),
    .Q(\rf.registers[19][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8869_ (.CLK(clk),
    .D(_0029_),
    .Q(\rf.registers[19][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8870_ (.CLK(clk),
    .D(_0030_),
    .Q(\rf.registers[19][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8871_ (.CLK(clk),
    .D(_0031_),
    .Q(\rf.registers[19][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8872_ (.CLK(clk),
    .D(_0032_),
    .Q(\rf.registers[19][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8873_ (.CLK(clk),
    .D(_0033_),
    .Q(\rf.registers[19][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8874_ (.CLK(clk),
    .D(_0034_),
    .Q(\rf.registers[19][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8875_ (.CLK(clk),
    .D(_0035_),
    .Q(\rf.registers[19][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8876_ (.CLK(clk),
    .D(_0036_),
    .Q(\rf.registers[19][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8877_ (.CLK(clk),
    .D(_0037_),
    .Q(\rf.registers[19][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8878_ (.CLK(clk),
    .D(_0038_),
    .Q(\rf.registers[19][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8879_ (.CLK(clk),
    .D(_0039_),
    .Q(\rf.registers[19][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8880_ (.CLK(clk),
    .D(_0040_),
    .Q(\rf.registers[19][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8881_ (.CLK(clk),
    .D(_0041_),
    .Q(\rf.registers[19][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8882_ (.CLK(clk),
    .D(_0042_),
    .Q(\rf.registers[19][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8883_ (.CLK(clk),
    .D(_0043_),
    .Q(\rf.registers[19][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8884_ (.CLK(clk),
    .D(_0044_),
    .Q(\rf.registers[19][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8885_ (.CLK(clk),
    .D(_0045_),
    .Q(\rf.registers[19][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8886_ (.CLK(clk),
    .D(_0046_),
    .Q(\rf.registers[19][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8887_ (.CLK(clk),
    .D(_0047_),
    .Q(\rf.registers[19][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8888_ (.CLK(clk),
    .D(_0048_),
    .Q(\rf.registers[19][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8889_ (.CLK(clk),
    .D(_0049_),
    .Q(\rf.registers[19][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8890_ (.CLK(clk),
    .D(_0050_),
    .Q(\rf.registers[19][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8891_ (.CLK(clk),
    .D(_0051_),
    .Q(\rf.registers[19][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8892_ (.CLK(clk),
    .D(_0052_),
    .Q(\rf.registers[19][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8893_ (.CLK(clk),
    .D(_0053_),
    .Q(\rf.registers[19][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8894_ (.CLK(clk),
    .D(_0054_),
    .Q(\rf.registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8895_ (.CLK(clk),
    .D(_0055_),
    .Q(\rf.registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8896_ (.CLK(clk),
    .D(_0056_),
    .Q(\rf.registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8897_ (.CLK(clk),
    .D(_0057_),
    .Q(\rf.registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8898_ (.CLK(clk),
    .D(_0058_),
    .Q(\rf.registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8899_ (.CLK(clk),
    .D(_0059_),
    .Q(\rf.registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8900_ (.CLK(clk),
    .D(_0060_),
    .Q(\rf.registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8901_ (.CLK(clk),
    .D(_0061_),
    .Q(\rf.registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8902_ (.CLK(clk),
    .D(_0062_),
    .Q(\rf.registers[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8903_ (.CLK(clk),
    .D(_0063_),
    .Q(\rf.registers[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8904_ (.CLK(clk),
    .D(_0064_),
    .Q(\rf.registers[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8905_ (.CLK(clk),
    .D(_0065_),
    .Q(\rf.registers[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8906_ (.CLK(clk),
    .D(_0066_),
    .Q(\rf.registers[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8907_ (.CLK(clk),
    .D(_0067_),
    .Q(\rf.registers[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8908_ (.CLK(clk),
    .D(_0068_),
    .Q(\rf.registers[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8909_ (.CLK(clk),
    .D(_0069_),
    .Q(\rf.registers[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8910_ (.CLK(clk),
    .D(_0070_),
    .Q(\rf.registers[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8911_ (.CLK(clk),
    .D(_0071_),
    .Q(\rf.registers[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8912_ (.CLK(clk),
    .D(_0072_),
    .Q(\rf.registers[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8913_ (.CLK(clk),
    .D(_0073_),
    .Q(\rf.registers[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8914_ (.CLK(clk),
    .D(_0074_),
    .Q(\rf.registers[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8915_ (.CLK(clk),
    .D(_0075_),
    .Q(\rf.registers[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8916_ (.CLK(clk),
    .D(_0076_),
    .Q(\rf.registers[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8917_ (.CLK(clk),
    .D(_0077_),
    .Q(\rf.registers[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8918_ (.CLK(clk),
    .D(_0078_),
    .Q(\rf.registers[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8919_ (.CLK(clk),
    .D(_0079_),
    .Q(\rf.registers[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8920_ (.CLK(clk),
    .D(_0080_),
    .Q(\rf.registers[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8921_ (.CLK(clk),
    .D(_0081_),
    .Q(\rf.registers[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8922_ (.CLK(clk),
    .D(_0082_),
    .Q(\rf.registers[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8923_ (.CLK(clk),
    .D(_0083_),
    .Q(\rf.registers[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8924_ (.CLK(clk),
    .D(_0084_),
    .Q(\rf.registers[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8925_ (.CLK(clk),
    .D(_0085_),
    .Q(\rf.registers[3][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8926_ (.CLK(clk),
    .D(_0086_),
    .Q(\rf.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8927_ (.CLK(clk),
    .D(_0087_),
    .Q(\rf.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8928_ (.CLK(clk),
    .D(_0088_),
    .Q(\rf.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8929_ (.CLK(clk),
    .D(_0089_),
    .Q(\rf.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8930_ (.CLK(clk),
    .D(_0090_),
    .Q(\rf.registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8931_ (.CLK(clk),
    .D(_0091_),
    .Q(\rf.registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8932_ (.CLK(clk),
    .D(_0092_),
    .Q(\rf.registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8933_ (.CLK(clk),
    .D(_0093_),
    .Q(\rf.registers[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8934_ (.CLK(clk),
    .D(_0094_),
    .Q(\rf.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8935_ (.CLK(clk),
    .D(_0095_),
    .Q(\rf.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8936_ (.CLK(clk),
    .D(_0096_),
    .Q(\rf.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8937_ (.CLK(clk),
    .D(_0097_),
    .Q(\rf.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8938_ (.CLK(clk),
    .D(_0098_),
    .Q(\rf.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8939_ (.CLK(clk),
    .D(_0099_),
    .Q(\rf.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8940_ (.CLK(clk),
    .D(_0100_),
    .Q(\rf.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8941_ (.CLK(clk),
    .D(_0101_),
    .Q(\rf.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8942_ (.CLK(clk),
    .D(_0102_),
    .Q(\rf.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8943_ (.CLK(clk),
    .D(_0103_),
    .Q(\rf.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8944_ (.CLK(clk),
    .D(_0104_),
    .Q(\rf.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8945_ (.CLK(clk),
    .D(_0105_),
    .Q(\rf.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8946_ (.CLK(clk),
    .D(_0106_),
    .Q(\rf.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8947_ (.CLK(clk),
    .D(_0107_),
    .Q(\rf.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8948_ (.CLK(clk),
    .D(_0108_),
    .Q(\rf.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8949_ (.CLK(clk),
    .D(_0109_),
    .Q(\rf.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8950_ (.CLK(clk),
    .D(_0110_),
    .Q(\rf.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8951_ (.CLK(clk),
    .D(_0111_),
    .Q(\rf.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8952_ (.CLK(clk),
    .D(_0112_),
    .Q(\rf.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8953_ (.CLK(clk),
    .D(_0113_),
    .Q(\rf.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8954_ (.CLK(clk),
    .D(_0114_),
    .Q(\rf.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8955_ (.CLK(clk),
    .D(_0115_),
    .Q(\rf.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8956_ (.CLK(clk),
    .D(_0116_),
    .Q(\rf.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8957_ (.CLK(clk),
    .D(_0117_),
    .Q(\rf.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8958_ (.CLK(clk),
    .D(_0118_),
    .Q(\rf.registers[29][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8959_ (.CLK(clk),
    .D(_0119_),
    .Q(\rf.registers[29][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8960_ (.CLK(clk),
    .D(_0120_),
    .Q(\rf.registers[29][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8961_ (.CLK(clk),
    .D(_0121_),
    .Q(\rf.registers[29][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8962_ (.CLK(clk),
    .D(_0122_),
    .Q(\rf.registers[29][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8963_ (.CLK(clk),
    .D(_0123_),
    .Q(\rf.registers[29][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8964_ (.CLK(clk),
    .D(_0124_),
    .Q(\rf.registers[29][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8965_ (.CLK(clk),
    .D(_0125_),
    .Q(\rf.registers[29][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8966_ (.CLK(clk),
    .D(_0126_),
    .Q(\rf.registers[29][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8967_ (.CLK(clk),
    .D(_0127_),
    .Q(\rf.registers[29][9] ));
 sky130_fd_sc_hd__dfxtp_2 _8968_ (.CLK(clk),
    .D(_0128_),
    .Q(\rf.registers[29][10] ));
 sky130_fd_sc_hd__dfxtp_2 _8969_ (.CLK(clk),
    .D(_0129_),
    .Q(\rf.registers[29][11] ));
 sky130_fd_sc_hd__dfxtp_2 _8970_ (.CLK(clk),
    .D(_0130_),
    .Q(\rf.registers[29][12] ));
 sky130_fd_sc_hd__dfxtp_2 _8971_ (.CLK(clk),
    .D(_0131_),
    .Q(\rf.registers[29][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8972_ (.CLK(clk),
    .D(_0132_),
    .Q(\rf.registers[29][14] ));
 sky130_fd_sc_hd__dfxtp_2 _8973_ (.CLK(clk),
    .D(_0133_),
    .Q(\rf.registers[29][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8974_ (.CLK(clk),
    .D(_0134_),
    .Q(\rf.registers[29][16] ));
 sky130_fd_sc_hd__dfxtp_2 _8975_ (.CLK(clk),
    .D(_0135_),
    .Q(\rf.registers[29][17] ));
 sky130_fd_sc_hd__dfxtp_2 _8976_ (.CLK(clk),
    .D(_0136_),
    .Q(\rf.registers[29][18] ));
 sky130_fd_sc_hd__dfxtp_2 _8977_ (.CLK(clk),
    .D(_0137_),
    .Q(\rf.registers[29][19] ));
 sky130_fd_sc_hd__dfxtp_2 _8978_ (.CLK(clk),
    .D(_0138_),
    .Q(\rf.registers[29][20] ));
 sky130_fd_sc_hd__dfxtp_2 _8979_ (.CLK(clk),
    .D(_0139_),
    .Q(\rf.registers[29][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8980_ (.CLK(clk),
    .D(_0140_),
    .Q(\rf.registers[29][22] ));
 sky130_fd_sc_hd__dfxtp_2 _8981_ (.CLK(clk),
    .D(_0141_),
    .Q(\rf.registers[29][23] ));
 sky130_fd_sc_hd__dfxtp_2 _8982_ (.CLK(clk),
    .D(_0142_),
    .Q(\rf.registers[29][24] ));
 sky130_fd_sc_hd__dfxtp_2 _8983_ (.CLK(clk),
    .D(_0143_),
    .Q(\rf.registers[29][25] ));
 sky130_fd_sc_hd__dfxtp_2 _8984_ (.CLK(clk),
    .D(_0144_),
    .Q(\rf.registers[29][26] ));
 sky130_fd_sc_hd__dfxtp_2 _8985_ (.CLK(clk),
    .D(_0145_),
    .Q(\rf.registers[29][27] ));
 sky130_fd_sc_hd__dfxtp_2 _8986_ (.CLK(clk),
    .D(_0146_),
    .Q(\rf.registers[29][28] ));
 sky130_fd_sc_hd__dfxtp_2 _8987_ (.CLK(clk),
    .D(_0147_),
    .Q(\rf.registers[29][29] ));
 sky130_fd_sc_hd__dfxtp_2 _8988_ (.CLK(clk),
    .D(_0148_),
    .Q(\rf.registers[29][30] ));
 sky130_fd_sc_hd__dfxtp_2 _8989_ (.CLK(clk),
    .D(_0149_),
    .Q(\rf.registers[29][31] ));
 sky130_fd_sc_hd__dfxtp_2 _8990_ (.CLK(clk),
    .D(_0150_),
    .Q(\rf.registers[31][0] ));
 sky130_fd_sc_hd__dfxtp_2 _8991_ (.CLK(clk),
    .D(_0151_),
    .Q(\rf.registers[31][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8992_ (.CLK(clk),
    .D(_0152_),
    .Q(\rf.registers[31][2] ));
 sky130_fd_sc_hd__dfxtp_2 _8993_ (.CLK(clk),
    .D(_0153_),
    .Q(\rf.registers[31][3] ));
 sky130_fd_sc_hd__dfxtp_2 _8994_ (.CLK(clk),
    .D(_0154_),
    .Q(\rf.registers[31][4] ));
 sky130_fd_sc_hd__dfxtp_2 _8995_ (.CLK(clk),
    .D(_0155_),
    .Q(\rf.registers[31][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8996_ (.CLK(clk),
    .D(_0156_),
    .Q(\rf.registers[31][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8997_ (.CLK(clk),
    .D(_0157_),
    .Q(\rf.registers[31][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8998_ (.CLK(clk),
    .D(_0158_),
    .Q(\rf.registers[31][8] ));
 sky130_fd_sc_hd__dfxtp_2 _8999_ (.CLK(clk),
    .D(_0159_),
    .Q(\rf.registers[31][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9000_ (.CLK(clk),
    .D(_0160_),
    .Q(\rf.registers[31][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9001_ (.CLK(clk),
    .D(_0161_),
    .Q(\rf.registers[31][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9002_ (.CLK(clk),
    .D(_0162_),
    .Q(\rf.registers[31][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9003_ (.CLK(clk),
    .D(_0163_),
    .Q(\rf.registers[31][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9004_ (.CLK(clk),
    .D(_0164_),
    .Q(\rf.registers[31][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9005_ (.CLK(clk),
    .D(_0165_),
    .Q(\rf.registers[31][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9006_ (.CLK(clk),
    .D(_0166_),
    .Q(\rf.registers[31][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9007_ (.CLK(clk),
    .D(_0167_),
    .Q(\rf.registers[31][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9008_ (.CLK(clk),
    .D(_0168_),
    .Q(\rf.registers[31][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9009_ (.CLK(clk),
    .D(_0169_),
    .Q(\rf.registers[31][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9010_ (.CLK(clk),
    .D(_0170_),
    .Q(\rf.registers[31][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9011_ (.CLK(clk),
    .D(_0171_),
    .Q(\rf.registers[31][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9012_ (.CLK(clk),
    .D(_0172_),
    .Q(\rf.registers[31][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9013_ (.CLK(clk),
    .D(_0173_),
    .Q(\rf.registers[31][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9014_ (.CLK(clk),
    .D(_0174_),
    .Q(\rf.registers[31][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9015_ (.CLK(clk),
    .D(_0175_),
    .Q(\rf.registers[31][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9016_ (.CLK(clk),
    .D(_0176_),
    .Q(\rf.registers[31][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9017_ (.CLK(clk),
    .D(_0177_),
    .Q(\rf.registers[31][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9018_ (.CLK(clk),
    .D(_0178_),
    .Q(\rf.registers[31][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9019_ (.CLK(clk),
    .D(_0179_),
    .Q(\rf.registers[31][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9020_ (.CLK(clk),
    .D(_0180_),
    .Q(\rf.registers[31][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9021_ (.CLK(clk),
    .D(_0181_),
    .Q(\rf.registers[31][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9022_ (.CLK(clk),
    .D(_0182_),
    .Q(\rf.registers[26][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9023_ (.CLK(clk),
    .D(_0183_),
    .Q(\rf.registers[26][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9024_ (.CLK(clk),
    .D(_0184_),
    .Q(\rf.registers[26][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9025_ (.CLK(clk),
    .D(_0185_),
    .Q(\rf.registers[26][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9026_ (.CLK(clk),
    .D(_0186_),
    .Q(\rf.registers[26][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9027_ (.CLK(clk),
    .D(_0187_),
    .Q(\rf.registers[26][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9028_ (.CLK(clk),
    .D(_0188_),
    .Q(\rf.registers[26][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9029_ (.CLK(clk),
    .D(_0189_),
    .Q(\rf.registers[26][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9030_ (.CLK(clk),
    .D(_0190_),
    .Q(\rf.registers[26][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9031_ (.CLK(clk),
    .D(_0191_),
    .Q(\rf.registers[26][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9032_ (.CLK(clk),
    .D(_0192_),
    .Q(\rf.registers[26][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9033_ (.CLK(clk),
    .D(_0193_),
    .Q(\rf.registers[26][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9034_ (.CLK(clk),
    .D(_0194_),
    .Q(\rf.registers[26][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9035_ (.CLK(clk),
    .D(_0195_),
    .Q(\rf.registers[26][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9036_ (.CLK(clk),
    .D(_0196_),
    .Q(\rf.registers[26][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9037_ (.CLK(clk),
    .D(_0197_),
    .Q(\rf.registers[26][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9038_ (.CLK(clk),
    .D(_0198_),
    .Q(\rf.registers[26][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9039_ (.CLK(clk),
    .D(_0199_),
    .Q(\rf.registers[26][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9040_ (.CLK(clk),
    .D(_0200_),
    .Q(\rf.registers[26][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9041_ (.CLK(clk),
    .D(_0201_),
    .Q(\rf.registers[26][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9042_ (.CLK(clk),
    .D(_0202_),
    .Q(\rf.registers[26][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9043_ (.CLK(clk),
    .D(_0203_),
    .Q(\rf.registers[26][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9044_ (.CLK(clk),
    .D(_0204_),
    .Q(\rf.registers[26][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9045_ (.CLK(clk),
    .D(_0205_),
    .Q(\rf.registers[26][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9046_ (.CLK(clk),
    .D(_0206_),
    .Q(\rf.registers[26][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9047_ (.CLK(clk),
    .D(_0207_),
    .Q(\rf.registers[26][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9048_ (.CLK(clk),
    .D(_0208_),
    .Q(\rf.registers[26][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9049_ (.CLK(clk),
    .D(_0209_),
    .Q(\rf.registers[26][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9050_ (.CLK(clk),
    .D(_0210_),
    .Q(\rf.registers[26][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9051_ (.CLK(clk),
    .D(_0211_),
    .Q(\rf.registers[26][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9052_ (.CLK(clk),
    .D(_0212_),
    .Q(\rf.registers[26][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9053_ (.CLK(clk),
    .D(_0213_),
    .Q(\rf.registers[26][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9054_ (.CLK(clk),
    .D(_0214_),
    .Q(\rf.registers[25][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9055_ (.CLK(clk),
    .D(_0215_),
    .Q(\rf.registers[25][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9056_ (.CLK(clk),
    .D(_0216_),
    .Q(\rf.registers[25][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9057_ (.CLK(clk),
    .D(_0217_),
    .Q(\rf.registers[25][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9058_ (.CLK(clk),
    .D(_0218_),
    .Q(\rf.registers[25][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9059_ (.CLK(clk),
    .D(_0219_),
    .Q(\rf.registers[25][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9060_ (.CLK(clk),
    .D(_0220_),
    .Q(\rf.registers[25][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9061_ (.CLK(clk),
    .D(_0221_),
    .Q(\rf.registers[25][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9062_ (.CLK(clk),
    .D(_0222_),
    .Q(\rf.registers[25][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9063_ (.CLK(clk),
    .D(_0223_),
    .Q(\rf.registers[25][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9064_ (.CLK(clk),
    .D(_0224_),
    .Q(\rf.registers[25][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9065_ (.CLK(clk),
    .D(_0225_),
    .Q(\rf.registers[25][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9066_ (.CLK(clk),
    .D(_0226_),
    .Q(\rf.registers[25][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9067_ (.CLK(clk),
    .D(_0227_),
    .Q(\rf.registers[25][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9068_ (.CLK(clk),
    .D(_0228_),
    .Q(\rf.registers[25][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9069_ (.CLK(clk),
    .D(_0229_),
    .Q(\rf.registers[25][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9070_ (.CLK(clk),
    .D(_0230_),
    .Q(\rf.registers[25][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9071_ (.CLK(clk),
    .D(_0231_),
    .Q(\rf.registers[25][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9072_ (.CLK(clk),
    .D(_0232_),
    .Q(\rf.registers[25][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9073_ (.CLK(clk),
    .D(_0233_),
    .Q(\rf.registers[25][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9074_ (.CLK(clk),
    .D(_0234_),
    .Q(\rf.registers[25][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9075_ (.CLK(clk),
    .D(_0235_),
    .Q(\rf.registers[25][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9076_ (.CLK(clk),
    .D(_0236_),
    .Q(\rf.registers[25][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9077_ (.CLK(clk),
    .D(_0237_),
    .Q(\rf.registers[25][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9078_ (.CLK(clk),
    .D(_0238_),
    .Q(\rf.registers[25][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9079_ (.CLK(clk),
    .D(_0239_),
    .Q(\rf.registers[25][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9080_ (.CLK(clk),
    .D(_0240_),
    .Q(\rf.registers[25][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9081_ (.CLK(clk),
    .D(_0241_),
    .Q(\rf.registers[25][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9082_ (.CLK(clk),
    .D(_0242_),
    .Q(\rf.registers[25][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9083_ (.CLK(clk),
    .D(_0243_),
    .Q(\rf.registers[25][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9084_ (.CLK(clk),
    .D(_0244_),
    .Q(\rf.registers[25][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9085_ (.CLK(clk),
    .D(_0245_),
    .Q(\rf.registers[25][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9086_ (.CLK(clk),
    .D(_0246_),
    .Q(\rf.registers[27][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9087_ (.CLK(clk),
    .D(_0247_),
    .Q(\rf.registers[27][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9088_ (.CLK(clk),
    .D(_0248_),
    .Q(\rf.registers[27][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9089_ (.CLK(clk),
    .D(_0249_),
    .Q(\rf.registers[27][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9090_ (.CLK(clk),
    .D(_0250_),
    .Q(\rf.registers[27][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9091_ (.CLK(clk),
    .D(_0251_),
    .Q(\rf.registers[27][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9092_ (.CLK(clk),
    .D(_0252_),
    .Q(\rf.registers[27][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9093_ (.CLK(clk),
    .D(_0253_),
    .Q(\rf.registers[27][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9094_ (.CLK(clk),
    .D(_0254_),
    .Q(\rf.registers[27][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9095_ (.CLK(clk),
    .D(_0255_),
    .Q(\rf.registers[27][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9096_ (.CLK(clk),
    .D(_0256_),
    .Q(\rf.registers[27][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9097_ (.CLK(clk),
    .D(_0257_),
    .Q(\rf.registers[27][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9098_ (.CLK(clk),
    .D(_0258_),
    .Q(\rf.registers[27][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9099_ (.CLK(clk),
    .D(_0259_),
    .Q(\rf.registers[27][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9100_ (.CLK(clk),
    .D(_0260_),
    .Q(\rf.registers[27][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9101_ (.CLK(clk),
    .D(_0261_),
    .Q(\rf.registers[27][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9102_ (.CLK(clk),
    .D(_0262_),
    .Q(\rf.registers[27][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9103_ (.CLK(clk),
    .D(_0263_),
    .Q(\rf.registers[27][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9104_ (.CLK(clk),
    .D(_0264_),
    .Q(\rf.registers[27][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9105_ (.CLK(clk),
    .D(_0265_),
    .Q(\rf.registers[27][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9106_ (.CLK(clk),
    .D(_0266_),
    .Q(\rf.registers[27][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9107_ (.CLK(clk),
    .D(_0267_),
    .Q(\rf.registers[27][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9108_ (.CLK(clk),
    .D(_0268_),
    .Q(\rf.registers[27][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9109_ (.CLK(clk),
    .D(_0269_),
    .Q(\rf.registers[27][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9110_ (.CLK(clk),
    .D(_0270_),
    .Q(\rf.registers[27][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9111_ (.CLK(clk),
    .D(_0271_),
    .Q(\rf.registers[27][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9112_ (.CLK(clk),
    .D(_0272_),
    .Q(\rf.registers[27][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9113_ (.CLK(clk),
    .D(_0273_),
    .Q(\rf.registers[27][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9114_ (.CLK(clk),
    .D(_0274_),
    .Q(\rf.registers[27][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9115_ (.CLK(clk),
    .D(_0275_),
    .Q(\rf.registers[27][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9116_ (.CLK(clk),
    .D(_0276_),
    .Q(\rf.registers[27][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9117_ (.CLK(clk),
    .D(_0277_),
    .Q(\rf.registers[27][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9118_ (.CLK(clk),
    .D(_0278_),
    .Q(\rf.registers[28][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9119_ (.CLK(clk),
    .D(_0279_),
    .Q(\rf.registers[28][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9120_ (.CLK(clk),
    .D(_0280_),
    .Q(\rf.registers[28][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9121_ (.CLK(clk),
    .D(_0281_),
    .Q(\rf.registers[28][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9122_ (.CLK(clk),
    .D(_0282_),
    .Q(\rf.registers[28][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9123_ (.CLK(clk),
    .D(_0283_),
    .Q(\rf.registers[28][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9124_ (.CLK(clk),
    .D(_0284_),
    .Q(\rf.registers[28][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9125_ (.CLK(clk),
    .D(_0285_),
    .Q(\rf.registers[28][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9126_ (.CLK(clk),
    .D(_0286_),
    .Q(\rf.registers[28][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9127_ (.CLK(clk),
    .D(_0287_),
    .Q(\rf.registers[28][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9128_ (.CLK(clk),
    .D(_0288_),
    .Q(\rf.registers[28][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9129_ (.CLK(clk),
    .D(_0289_),
    .Q(\rf.registers[28][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9130_ (.CLK(clk),
    .D(_0290_),
    .Q(\rf.registers[28][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9131_ (.CLK(clk),
    .D(_0291_),
    .Q(\rf.registers[28][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9132_ (.CLK(clk),
    .D(_0292_),
    .Q(\rf.registers[28][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9133_ (.CLK(clk),
    .D(_0293_),
    .Q(\rf.registers[28][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9134_ (.CLK(clk),
    .D(_0294_),
    .Q(\rf.registers[28][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9135_ (.CLK(clk),
    .D(_0295_),
    .Q(\rf.registers[28][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9136_ (.CLK(clk),
    .D(_0296_),
    .Q(\rf.registers[28][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9137_ (.CLK(clk),
    .D(_0297_),
    .Q(\rf.registers[28][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9138_ (.CLK(clk),
    .D(_0298_),
    .Q(\rf.registers[28][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9139_ (.CLK(clk),
    .D(_0299_),
    .Q(\rf.registers[28][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9140_ (.CLK(clk),
    .D(_0300_),
    .Q(\rf.registers[28][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9141_ (.CLK(clk),
    .D(_0301_),
    .Q(\rf.registers[28][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9142_ (.CLK(clk),
    .D(_0302_),
    .Q(\rf.registers[28][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9143_ (.CLK(clk),
    .D(_0303_),
    .Q(\rf.registers[28][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9144_ (.CLK(clk),
    .D(_0304_),
    .Q(\rf.registers[28][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9145_ (.CLK(clk),
    .D(_0305_),
    .Q(\rf.registers[28][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9146_ (.CLK(clk),
    .D(_0306_),
    .Q(\rf.registers[28][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9147_ (.CLK(clk),
    .D(_0307_),
    .Q(\rf.registers[28][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9148_ (.CLK(clk),
    .D(_0308_),
    .Q(\rf.registers[28][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9149_ (.CLK(clk),
    .D(_0309_),
    .Q(\rf.registers[28][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9150_ (.CLK(clk),
    .D(_0310_),
    .Q(\rf.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9151_ (.CLK(clk),
    .D(_0311_),
    .Q(\rf.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9152_ (.CLK(clk),
    .D(_0312_),
    .Q(\rf.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9153_ (.CLK(clk),
    .D(_0313_),
    .Q(\rf.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9154_ (.CLK(clk),
    .D(_0314_),
    .Q(\rf.registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9155_ (.CLK(clk),
    .D(_0315_),
    .Q(\rf.registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9156_ (.CLK(clk),
    .D(_0316_),
    .Q(\rf.registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9157_ (.CLK(clk),
    .D(_0317_),
    .Q(\rf.registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9158_ (.CLK(clk),
    .D(_0318_),
    .Q(\rf.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9159_ (.CLK(clk),
    .D(_0319_),
    .Q(\rf.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9160_ (.CLK(clk),
    .D(_0320_),
    .Q(\rf.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9161_ (.CLK(clk),
    .D(_0321_),
    .Q(\rf.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9162_ (.CLK(clk),
    .D(_0322_),
    .Q(\rf.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9163_ (.CLK(clk),
    .D(_0323_),
    .Q(\rf.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9164_ (.CLK(clk),
    .D(_0324_),
    .Q(\rf.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9165_ (.CLK(clk),
    .D(_0325_),
    .Q(\rf.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9166_ (.CLK(clk),
    .D(_0326_),
    .Q(\rf.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9167_ (.CLK(clk),
    .D(_0327_),
    .Q(\rf.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9168_ (.CLK(clk),
    .D(_0328_),
    .Q(\rf.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9169_ (.CLK(clk),
    .D(_0329_),
    .Q(\rf.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9170_ (.CLK(clk),
    .D(_0330_),
    .Q(\rf.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9171_ (.CLK(clk),
    .D(_0331_),
    .Q(\rf.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9172_ (.CLK(clk),
    .D(_0332_),
    .Q(\rf.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9173_ (.CLK(clk),
    .D(_0333_),
    .Q(\rf.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9174_ (.CLK(clk),
    .D(_0334_),
    .Q(\rf.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9175_ (.CLK(clk),
    .D(_0335_),
    .Q(\rf.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9176_ (.CLK(clk),
    .D(_0336_),
    .Q(\rf.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9177_ (.CLK(clk),
    .D(_0337_),
    .Q(\rf.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9178_ (.CLK(clk),
    .D(_0338_),
    .Q(\rf.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9179_ (.CLK(clk),
    .D(_0339_),
    .Q(\rf.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9180_ (.CLK(clk),
    .D(_0340_),
    .Q(\rf.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9181_ (.CLK(clk),
    .D(_0341_),
    .Q(\rf.registers[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9182_ (.CLK(clk),
    .D(_0342_),
    .Q(\rf.registers[30][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9183_ (.CLK(clk),
    .D(_0343_),
    .Q(\rf.registers[30][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9184_ (.CLK(clk),
    .D(_0344_),
    .Q(\rf.registers[30][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9185_ (.CLK(clk),
    .D(_0345_),
    .Q(\rf.registers[30][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9186_ (.CLK(clk),
    .D(_0346_),
    .Q(\rf.registers[30][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9187_ (.CLK(clk),
    .D(_0347_),
    .Q(\rf.registers[30][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9188_ (.CLK(clk),
    .D(_0348_),
    .Q(\rf.registers[30][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9189_ (.CLK(clk),
    .D(_0349_),
    .Q(\rf.registers[30][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9190_ (.CLK(clk),
    .D(_0350_),
    .Q(\rf.registers[30][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9191_ (.CLK(clk),
    .D(_0351_),
    .Q(\rf.registers[30][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9192_ (.CLK(clk),
    .D(_0352_),
    .Q(\rf.registers[30][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9193_ (.CLK(clk),
    .D(_0353_),
    .Q(\rf.registers[30][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9194_ (.CLK(clk),
    .D(_0354_),
    .Q(\rf.registers[30][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9195_ (.CLK(clk),
    .D(_0355_),
    .Q(\rf.registers[30][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9196_ (.CLK(clk),
    .D(_0356_),
    .Q(\rf.registers[30][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9197_ (.CLK(clk),
    .D(_0357_),
    .Q(\rf.registers[30][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9198_ (.CLK(clk),
    .D(_0358_),
    .Q(\rf.registers[30][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9199_ (.CLK(clk),
    .D(_0359_),
    .Q(\rf.registers[30][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9200_ (.CLK(clk),
    .D(_0360_),
    .Q(\rf.registers[30][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9201_ (.CLK(clk),
    .D(_0361_),
    .Q(\rf.registers[30][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9202_ (.CLK(clk),
    .D(_0362_),
    .Q(\rf.registers[30][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9203_ (.CLK(clk),
    .D(_0363_),
    .Q(\rf.registers[30][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9204_ (.CLK(clk),
    .D(_0364_),
    .Q(\rf.registers[30][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9205_ (.CLK(clk),
    .D(_0365_),
    .Q(\rf.registers[30][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9206_ (.CLK(clk),
    .D(_0366_),
    .Q(\rf.registers[30][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9207_ (.CLK(clk),
    .D(_0367_),
    .Q(\rf.registers[30][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9208_ (.CLK(clk),
    .D(_0368_),
    .Q(\rf.registers[30][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9209_ (.CLK(clk),
    .D(_0369_),
    .Q(\rf.registers[30][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9210_ (.CLK(clk),
    .D(_0370_),
    .Q(\rf.registers[30][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9211_ (.CLK(clk),
    .D(_0371_),
    .Q(\rf.registers[30][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9212_ (.CLK(clk),
    .D(_0372_),
    .Q(\rf.registers[30][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9213_ (.CLK(clk),
    .D(_0373_),
    .Q(\rf.registers[30][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9214_ (.CLK(clk),
    .D(_0374_),
    .Q(\rf.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9215_ (.CLK(clk),
    .D(_0375_),
    .Q(\rf.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9216_ (.CLK(clk),
    .D(_0376_),
    .Q(\rf.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9217_ (.CLK(clk),
    .D(_0377_),
    .Q(\rf.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9218_ (.CLK(clk),
    .D(_0378_),
    .Q(\rf.registers[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9219_ (.CLK(clk),
    .D(_0379_),
    .Q(\rf.registers[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9220_ (.CLK(clk),
    .D(_0380_),
    .Q(\rf.registers[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9221_ (.CLK(clk),
    .D(_0381_),
    .Q(\rf.registers[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9222_ (.CLK(clk),
    .D(_0382_),
    .Q(\rf.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9223_ (.CLK(clk),
    .D(_0383_),
    .Q(\rf.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9224_ (.CLK(clk),
    .D(_0384_),
    .Q(\rf.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9225_ (.CLK(clk),
    .D(_0385_),
    .Q(\rf.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9226_ (.CLK(clk),
    .D(_0386_),
    .Q(\rf.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9227_ (.CLK(clk),
    .D(_0387_),
    .Q(\rf.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9228_ (.CLK(clk),
    .D(_0388_),
    .Q(\rf.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9229_ (.CLK(clk),
    .D(_0389_),
    .Q(\rf.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9230_ (.CLK(clk),
    .D(_0390_),
    .Q(\rf.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9231_ (.CLK(clk),
    .D(_0391_),
    .Q(\rf.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9232_ (.CLK(clk),
    .D(_0392_),
    .Q(\rf.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9233_ (.CLK(clk),
    .D(_0393_),
    .Q(\rf.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9234_ (.CLK(clk),
    .D(_0394_),
    .Q(\rf.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9235_ (.CLK(clk),
    .D(_0395_),
    .Q(\rf.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9236_ (.CLK(clk),
    .D(_0396_),
    .Q(\rf.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9237_ (.CLK(clk),
    .D(_0397_),
    .Q(\rf.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9238_ (.CLK(clk),
    .D(_0398_),
    .Q(\rf.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9239_ (.CLK(clk),
    .D(_0399_),
    .Q(\rf.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9240_ (.CLK(clk),
    .D(_0400_),
    .Q(\rf.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9241_ (.CLK(clk),
    .D(_0401_),
    .Q(\rf.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9242_ (.CLK(clk),
    .D(_0402_),
    .Q(\rf.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9243_ (.CLK(clk),
    .D(_0403_),
    .Q(\rf.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9244_ (.CLK(clk),
    .D(_0404_),
    .Q(\rf.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9245_ (.CLK(clk),
    .D(_0405_),
    .Q(\rf.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9246_ (.CLK(clk),
    .D(_0406_),
    .Q(\rf.registers[23][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9247_ (.CLK(clk),
    .D(_0407_),
    .Q(\rf.registers[23][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9248_ (.CLK(clk),
    .D(_0408_),
    .Q(\rf.registers[23][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9249_ (.CLK(clk),
    .D(_0409_),
    .Q(\rf.registers[23][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9250_ (.CLK(clk),
    .D(_0410_),
    .Q(\rf.registers[23][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9251_ (.CLK(clk),
    .D(_0411_),
    .Q(\rf.registers[23][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9252_ (.CLK(clk),
    .D(_0412_),
    .Q(\rf.registers[23][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9253_ (.CLK(clk),
    .D(_0413_),
    .Q(\rf.registers[23][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9254_ (.CLK(clk),
    .D(_0414_),
    .Q(\rf.registers[23][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9255_ (.CLK(clk),
    .D(_0415_),
    .Q(\rf.registers[23][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9256_ (.CLK(clk),
    .D(_0416_),
    .Q(\rf.registers[23][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9257_ (.CLK(clk),
    .D(_0417_),
    .Q(\rf.registers[23][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9258_ (.CLK(clk),
    .D(_0418_),
    .Q(\rf.registers[23][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9259_ (.CLK(clk),
    .D(_0419_),
    .Q(\rf.registers[23][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9260_ (.CLK(clk),
    .D(_0420_),
    .Q(\rf.registers[23][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9261_ (.CLK(clk),
    .D(_0421_),
    .Q(\rf.registers[23][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9262_ (.CLK(clk),
    .D(_0422_),
    .Q(\rf.registers[23][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9263_ (.CLK(clk),
    .D(_0423_),
    .Q(\rf.registers[23][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9264_ (.CLK(clk),
    .D(_0424_),
    .Q(\rf.registers[23][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9265_ (.CLK(clk),
    .D(_0425_),
    .Q(\rf.registers[23][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9266_ (.CLK(clk),
    .D(_0426_),
    .Q(\rf.registers[23][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9267_ (.CLK(clk),
    .D(_0427_),
    .Q(\rf.registers[23][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9268_ (.CLK(clk),
    .D(_0428_),
    .Q(\rf.registers[23][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9269_ (.CLK(clk),
    .D(_0429_),
    .Q(\rf.registers[23][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9270_ (.CLK(clk),
    .D(_0430_),
    .Q(\rf.registers[23][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9271_ (.CLK(clk),
    .D(_0431_),
    .Q(\rf.registers[23][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9272_ (.CLK(clk),
    .D(_0432_),
    .Q(\rf.registers[23][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9273_ (.CLK(clk),
    .D(_0433_),
    .Q(\rf.registers[23][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9274_ (.CLK(clk),
    .D(_0434_),
    .Q(\rf.registers[23][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9275_ (.CLK(clk),
    .D(_0435_),
    .Q(\rf.registers[23][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9276_ (.CLK(clk),
    .D(_0436_),
    .Q(\rf.registers[23][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9277_ (.CLK(clk),
    .D(_0437_),
    .Q(\rf.registers[23][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9278_ (.CLK(clk),
    .D(_0438_),
    .Q(\rf.registers[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9279_ (.CLK(clk),
    .D(_0439_),
    .Q(\rf.registers[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9280_ (.CLK(clk),
    .D(_0440_),
    .Q(\rf.registers[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9281_ (.CLK(clk),
    .D(_0441_),
    .Q(\rf.registers[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9282_ (.CLK(clk),
    .D(_0442_),
    .Q(\rf.registers[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9283_ (.CLK(clk),
    .D(_0443_),
    .Q(\rf.registers[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9284_ (.CLK(clk),
    .D(_0444_),
    .Q(\rf.registers[18][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9285_ (.CLK(clk),
    .D(_0445_),
    .Q(\rf.registers[18][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9286_ (.CLK(clk),
    .D(_0446_),
    .Q(\rf.registers[18][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9287_ (.CLK(clk),
    .D(_0447_),
    .Q(\rf.registers[18][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9288_ (.CLK(clk),
    .D(_0448_),
    .Q(\rf.registers[18][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9289_ (.CLK(clk),
    .D(_0449_),
    .Q(\rf.registers[18][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9290_ (.CLK(clk),
    .D(_0450_),
    .Q(\rf.registers[18][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9291_ (.CLK(clk),
    .D(_0451_),
    .Q(\rf.registers[18][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9292_ (.CLK(clk),
    .D(_0452_),
    .Q(\rf.registers[18][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9293_ (.CLK(clk),
    .D(_0453_),
    .Q(\rf.registers[18][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9294_ (.CLK(clk),
    .D(_0454_),
    .Q(\rf.registers[18][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9295_ (.CLK(clk),
    .D(_0455_),
    .Q(\rf.registers[18][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9296_ (.CLK(clk),
    .D(_0456_),
    .Q(\rf.registers[18][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9297_ (.CLK(clk),
    .D(_0457_),
    .Q(\rf.registers[18][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9298_ (.CLK(clk),
    .D(_0458_),
    .Q(\rf.registers[18][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9299_ (.CLK(clk),
    .D(_0459_),
    .Q(\rf.registers[18][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9300_ (.CLK(clk),
    .D(_0460_),
    .Q(\rf.registers[18][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9301_ (.CLK(clk),
    .D(_0461_),
    .Q(\rf.registers[18][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9302_ (.CLK(clk),
    .D(_0462_),
    .Q(\rf.registers[18][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9303_ (.CLK(clk),
    .D(_0463_),
    .Q(\rf.registers[18][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9304_ (.CLK(clk),
    .D(_0464_),
    .Q(\rf.registers[18][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9305_ (.CLK(clk),
    .D(_0465_),
    .Q(\rf.registers[18][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9306_ (.CLK(clk),
    .D(_0466_),
    .Q(\rf.registers[18][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9307_ (.CLK(clk),
    .D(_0467_),
    .Q(\rf.registers[18][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9308_ (.CLK(clk),
    .D(_0468_),
    .Q(\rf.registers[18][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9309_ (.CLK(clk),
    .D(_0469_),
    .Q(\rf.registers[18][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9310_ (.CLK(clk),
    .D(_0470_),
    .Q(\rf.registers[21][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9311_ (.CLK(clk),
    .D(_0471_),
    .Q(\rf.registers[21][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9312_ (.CLK(clk),
    .D(_0472_),
    .Q(\rf.registers[21][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9313_ (.CLK(clk),
    .D(_0473_),
    .Q(\rf.registers[21][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9314_ (.CLK(clk),
    .D(_0474_),
    .Q(\rf.registers[21][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9315_ (.CLK(clk),
    .D(_0475_),
    .Q(\rf.registers[21][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9316_ (.CLK(clk),
    .D(_0476_),
    .Q(\rf.registers[21][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9317_ (.CLK(clk),
    .D(_0477_),
    .Q(\rf.registers[21][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9318_ (.CLK(clk),
    .D(_0478_),
    .Q(\rf.registers[21][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9319_ (.CLK(clk),
    .D(_0479_),
    .Q(\rf.registers[21][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9320_ (.CLK(clk),
    .D(_0480_),
    .Q(\rf.registers[21][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9321_ (.CLK(clk),
    .D(_0481_),
    .Q(\rf.registers[21][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9322_ (.CLK(clk),
    .D(_0482_),
    .Q(\rf.registers[21][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9323_ (.CLK(clk),
    .D(_0483_),
    .Q(\rf.registers[21][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9324_ (.CLK(clk),
    .D(_0484_),
    .Q(\rf.registers[21][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9325_ (.CLK(clk),
    .D(_0485_),
    .Q(\rf.registers[21][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9326_ (.CLK(clk),
    .D(_0486_),
    .Q(\rf.registers[21][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9327_ (.CLK(clk),
    .D(_0487_),
    .Q(\rf.registers[21][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9328_ (.CLK(clk),
    .D(_0488_),
    .Q(\rf.registers[21][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9329_ (.CLK(clk),
    .D(_0489_),
    .Q(\rf.registers[21][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9330_ (.CLK(clk),
    .D(_0490_),
    .Q(\rf.registers[21][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9331_ (.CLK(clk),
    .D(_0491_),
    .Q(\rf.registers[21][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9332_ (.CLK(clk),
    .D(_0492_),
    .Q(\rf.registers[21][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9333_ (.CLK(clk),
    .D(_0493_),
    .Q(\rf.registers[21][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9334_ (.CLK(clk),
    .D(_0494_),
    .Q(\rf.registers[21][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9335_ (.CLK(clk),
    .D(_0495_),
    .Q(\rf.registers[21][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9336_ (.CLK(clk),
    .D(_0496_),
    .Q(\rf.registers[21][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9337_ (.CLK(clk),
    .D(_0497_),
    .Q(\rf.registers[21][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9338_ (.CLK(clk),
    .D(_0498_),
    .Q(\rf.registers[21][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9339_ (.CLK(clk),
    .D(_0499_),
    .Q(\rf.registers[21][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9340_ (.CLK(clk),
    .D(_0500_),
    .Q(\rf.registers[21][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9341_ (.CLK(clk),
    .D(_0501_),
    .Q(\rf.registers[21][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9342_ (.CLK(clk),
    .D(_0502_),
    .Q(\rf.registers[20][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9343_ (.CLK(clk),
    .D(_0503_),
    .Q(\rf.registers[20][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9344_ (.CLK(clk),
    .D(_0504_),
    .Q(\rf.registers[20][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9345_ (.CLK(clk),
    .D(_0505_),
    .Q(\rf.registers[20][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9346_ (.CLK(clk),
    .D(_0506_),
    .Q(\rf.registers[20][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9347_ (.CLK(clk),
    .D(_0507_),
    .Q(\rf.registers[20][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9348_ (.CLK(clk),
    .D(_0508_),
    .Q(\rf.registers[20][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9349_ (.CLK(clk),
    .D(_0509_),
    .Q(\rf.registers[20][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9350_ (.CLK(clk),
    .D(_0510_),
    .Q(\rf.registers[20][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9351_ (.CLK(clk),
    .D(_0511_),
    .Q(\rf.registers[20][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9352_ (.CLK(clk),
    .D(_0512_),
    .Q(\rf.registers[20][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9353_ (.CLK(clk),
    .D(_0513_),
    .Q(\rf.registers[20][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9354_ (.CLK(clk),
    .D(_0514_),
    .Q(\rf.registers[20][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9355_ (.CLK(clk),
    .D(_0515_),
    .Q(\rf.registers[20][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9356_ (.CLK(clk),
    .D(_0516_),
    .Q(\rf.registers[20][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9357_ (.CLK(clk),
    .D(_0517_),
    .Q(\rf.registers[20][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9358_ (.CLK(clk),
    .D(_0518_),
    .Q(\rf.registers[20][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9359_ (.CLK(clk),
    .D(_0519_),
    .Q(\rf.registers[20][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9360_ (.CLK(clk),
    .D(_0520_),
    .Q(\rf.registers[20][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9361_ (.CLK(clk),
    .D(_0521_),
    .Q(\rf.registers[20][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9362_ (.CLK(clk),
    .D(_0522_),
    .Q(\rf.registers[20][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9363_ (.CLK(clk),
    .D(_0523_),
    .Q(\rf.registers[20][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9364_ (.CLK(clk),
    .D(_0524_),
    .Q(\rf.registers[20][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9365_ (.CLK(clk),
    .D(_0525_),
    .Q(\rf.registers[20][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9366_ (.CLK(clk),
    .D(_0526_),
    .Q(\rf.registers[20][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9367_ (.CLK(clk),
    .D(_0527_),
    .Q(\rf.registers[20][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9368_ (.CLK(clk),
    .D(_0528_),
    .Q(\rf.registers[20][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9369_ (.CLK(clk),
    .D(_0529_),
    .Q(\rf.registers[20][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9370_ (.CLK(clk),
    .D(_0530_),
    .Q(\rf.registers[20][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9371_ (.CLK(clk),
    .D(_0531_),
    .Q(\rf.registers[20][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9372_ (.CLK(clk),
    .D(_0532_),
    .Q(\rf.registers[20][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9373_ (.CLK(clk),
    .D(_0533_),
    .Q(\rf.registers[20][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9374_ (.CLK(clk),
    .D(_0534_),
    .Q(\rf.registers[24][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9375_ (.CLK(clk),
    .D(_0535_),
    .Q(\rf.registers[24][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9376_ (.CLK(clk),
    .D(_0536_),
    .Q(\rf.registers[24][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9377_ (.CLK(clk),
    .D(_0537_),
    .Q(\rf.registers[24][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9378_ (.CLK(clk),
    .D(_0538_),
    .Q(\rf.registers[24][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9379_ (.CLK(clk),
    .D(_0539_),
    .Q(\rf.registers[24][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9380_ (.CLK(clk),
    .D(_0540_),
    .Q(\rf.registers[24][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9381_ (.CLK(clk),
    .D(_0541_),
    .Q(\rf.registers[24][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9382_ (.CLK(clk),
    .D(_0542_),
    .Q(\rf.registers[24][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9383_ (.CLK(clk),
    .D(_0543_),
    .Q(\rf.registers[24][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9384_ (.CLK(clk),
    .D(_0544_),
    .Q(\rf.registers[24][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9385_ (.CLK(clk),
    .D(_0545_),
    .Q(\rf.registers[24][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9386_ (.CLK(clk),
    .D(_0546_),
    .Q(\rf.registers[24][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9387_ (.CLK(clk),
    .D(_0547_),
    .Q(\rf.registers[24][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9388_ (.CLK(clk),
    .D(_0548_),
    .Q(\rf.registers[24][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9389_ (.CLK(clk),
    .D(_0549_),
    .Q(\rf.registers[24][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9390_ (.CLK(clk),
    .D(_0550_),
    .Q(\rf.registers[24][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9391_ (.CLK(clk),
    .D(_0551_),
    .Q(\rf.registers[24][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9392_ (.CLK(clk),
    .D(_0552_),
    .Q(\rf.registers[24][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9393_ (.CLK(clk),
    .D(_0553_),
    .Q(\rf.registers[24][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9394_ (.CLK(clk),
    .D(_0554_),
    .Q(\rf.registers[24][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9395_ (.CLK(clk),
    .D(_0555_),
    .Q(\rf.registers[24][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9396_ (.CLK(clk),
    .D(_0556_),
    .Q(\rf.registers[24][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9397_ (.CLK(clk),
    .D(_0557_),
    .Q(\rf.registers[24][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9398_ (.CLK(clk),
    .D(_0558_),
    .Q(\rf.registers[24][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9399_ (.CLK(clk),
    .D(_0559_),
    .Q(\rf.registers[24][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9400_ (.CLK(clk),
    .D(_0560_),
    .Q(\rf.registers[24][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9401_ (.CLK(clk),
    .D(_0561_),
    .Q(\rf.registers[24][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9402_ (.CLK(clk),
    .D(_0562_),
    .Q(\rf.registers[24][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9403_ (.CLK(clk),
    .D(_0563_),
    .Q(\rf.registers[24][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9404_ (.CLK(clk),
    .D(_0564_),
    .Q(\rf.registers[24][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9405_ (.CLK(clk),
    .D(_0565_),
    .Q(\rf.registers[24][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9406_ (.CLK(clk),
    .D(_0566_),
    .Q(\rf.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9407_ (.CLK(clk),
    .D(_0567_),
    .Q(\rf.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9408_ (.CLK(clk),
    .D(_0568_),
    .Q(\rf.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9409_ (.CLK(clk),
    .D(_0569_),
    .Q(\rf.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9410_ (.CLK(clk),
    .D(_0570_),
    .Q(\rf.registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9411_ (.CLK(clk),
    .D(_0571_),
    .Q(\rf.registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9412_ (.CLK(clk),
    .D(_0572_),
    .Q(\rf.registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9413_ (.CLK(clk),
    .D(_0573_),
    .Q(\rf.registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9414_ (.CLK(clk),
    .D(_0574_),
    .Q(\rf.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9415_ (.CLK(clk),
    .D(_0575_),
    .Q(\rf.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9416_ (.CLK(clk),
    .D(_0576_),
    .Q(\rf.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9417_ (.CLK(clk),
    .D(_0577_),
    .Q(\rf.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9418_ (.CLK(clk),
    .D(_0578_),
    .Q(\rf.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9419_ (.CLK(clk),
    .D(_0579_),
    .Q(\rf.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9420_ (.CLK(clk),
    .D(_0580_),
    .Q(\rf.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9421_ (.CLK(clk),
    .D(_0581_),
    .Q(\rf.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9422_ (.CLK(clk),
    .D(_0582_),
    .Q(\rf.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9423_ (.CLK(clk),
    .D(_0583_),
    .Q(\rf.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9424_ (.CLK(clk),
    .D(_0584_),
    .Q(\rf.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9425_ (.CLK(clk),
    .D(_0585_),
    .Q(\rf.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9426_ (.CLK(clk),
    .D(_0586_),
    .Q(\rf.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9427_ (.CLK(clk),
    .D(_0587_),
    .Q(\rf.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9428_ (.CLK(clk),
    .D(_0588_),
    .Q(\rf.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9429_ (.CLK(clk),
    .D(_0589_),
    .Q(\rf.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9430_ (.CLK(clk),
    .D(_0590_),
    .Q(\rf.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9431_ (.CLK(clk),
    .D(_0591_),
    .Q(\rf.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9432_ (.CLK(clk),
    .D(_0592_),
    .Q(\rf.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9433_ (.CLK(clk),
    .D(_0593_),
    .Q(\rf.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9434_ (.CLK(clk),
    .D(_0594_),
    .Q(\rf.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9435_ (.CLK(clk),
    .D(_0595_),
    .Q(\rf.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9436_ (.CLK(clk),
    .D(_0596_),
    .Q(\rf.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9437_ (.CLK(clk),
    .D(_0597_),
    .Q(\rf.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9438_ (.CLK(clk),
    .D(_0598_),
    .Q(\rf.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9439_ (.CLK(clk),
    .D(_0599_),
    .Q(\rf.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9440_ (.CLK(clk),
    .D(_0600_),
    .Q(\rf.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9441_ (.CLK(clk),
    .D(_0601_),
    .Q(\rf.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9442_ (.CLK(clk),
    .D(_0602_),
    .Q(\rf.registers[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9443_ (.CLK(clk),
    .D(_0603_),
    .Q(\rf.registers[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9444_ (.CLK(clk),
    .D(_0604_),
    .Q(\rf.registers[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9445_ (.CLK(clk),
    .D(_0605_),
    .Q(\rf.registers[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9446_ (.CLK(clk),
    .D(_0606_),
    .Q(\rf.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9447_ (.CLK(clk),
    .D(_0607_),
    .Q(\rf.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9448_ (.CLK(clk),
    .D(_0608_),
    .Q(\rf.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9449_ (.CLK(clk),
    .D(_0609_),
    .Q(\rf.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9450_ (.CLK(clk),
    .D(_0610_),
    .Q(\rf.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9451_ (.CLK(clk),
    .D(_0611_),
    .Q(\rf.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9452_ (.CLK(clk),
    .D(_0612_),
    .Q(\rf.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9453_ (.CLK(clk),
    .D(_0613_),
    .Q(\rf.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9454_ (.CLK(clk),
    .D(_0614_),
    .Q(\rf.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9455_ (.CLK(clk),
    .D(_0615_),
    .Q(\rf.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9456_ (.CLK(clk),
    .D(_0616_),
    .Q(\rf.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9457_ (.CLK(clk),
    .D(_0617_),
    .Q(\rf.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9458_ (.CLK(clk),
    .D(_0618_),
    .Q(\rf.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9459_ (.CLK(clk),
    .D(_0619_),
    .Q(\rf.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9460_ (.CLK(clk),
    .D(_0620_),
    .Q(\rf.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9461_ (.CLK(clk),
    .D(_0621_),
    .Q(\rf.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9462_ (.CLK(clk),
    .D(_0622_),
    .Q(\rf.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9463_ (.CLK(clk),
    .D(_0623_),
    .Q(\rf.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9464_ (.CLK(clk),
    .D(_0624_),
    .Q(\rf.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9465_ (.CLK(clk),
    .D(_0625_),
    .Q(\rf.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9466_ (.CLK(clk),
    .D(_0626_),
    .Q(\rf.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9467_ (.CLK(clk),
    .D(_0627_),
    .Q(\rf.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9468_ (.CLK(clk),
    .D(_0628_),
    .Q(\rf.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9469_ (.CLK(clk),
    .D(_0629_),
    .Q(\rf.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9470_ (.CLK(clk),
    .D(_0630_),
    .Q(\rf.registers[16][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9471_ (.CLK(clk),
    .D(_0631_),
    .Q(\rf.registers[16][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9472_ (.CLK(clk),
    .D(_0632_),
    .Q(\rf.registers[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9473_ (.CLK(clk),
    .D(_0633_),
    .Q(\rf.registers[16][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9474_ (.CLK(clk),
    .D(_0634_),
    .Q(\rf.registers[16][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9475_ (.CLK(clk),
    .D(_0635_),
    .Q(\rf.registers[16][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9476_ (.CLK(clk),
    .D(_0636_),
    .Q(\rf.registers[16][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9477_ (.CLK(clk),
    .D(_0637_),
    .Q(\rf.registers[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9478_ (.CLK(clk),
    .D(_0638_),
    .Q(\rf.registers[16][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9479_ (.CLK(clk),
    .D(_0639_),
    .Q(\rf.registers[16][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9480_ (.CLK(clk),
    .D(_0640_),
    .Q(\rf.registers[16][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9481_ (.CLK(clk),
    .D(_0641_),
    .Q(\rf.registers[16][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9482_ (.CLK(clk),
    .D(_0642_),
    .Q(\rf.registers[16][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9483_ (.CLK(clk),
    .D(_0643_),
    .Q(\rf.registers[16][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9484_ (.CLK(clk),
    .D(_0644_),
    .Q(\rf.registers[16][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9485_ (.CLK(clk),
    .D(_0645_),
    .Q(\rf.registers[16][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9486_ (.CLK(clk),
    .D(_0646_),
    .Q(\rf.registers[16][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9487_ (.CLK(clk),
    .D(_0647_),
    .Q(\rf.registers[16][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9488_ (.CLK(clk),
    .D(_0648_),
    .Q(\rf.registers[16][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9489_ (.CLK(clk),
    .D(_0649_),
    .Q(\rf.registers[16][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9490_ (.CLK(clk),
    .D(_0650_),
    .Q(\rf.registers[16][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9491_ (.CLK(clk),
    .D(_0651_),
    .Q(\rf.registers[16][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9492_ (.CLK(clk),
    .D(_0652_),
    .Q(\rf.registers[16][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9493_ (.CLK(clk),
    .D(_0653_),
    .Q(\rf.registers[16][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9494_ (.CLK(clk),
    .D(_0654_),
    .Q(\rf.registers[16][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9495_ (.CLK(clk),
    .D(_0655_),
    .Q(\rf.registers[16][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9496_ (.CLK(clk),
    .D(_0656_),
    .Q(\rf.registers[16][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9497_ (.CLK(clk),
    .D(_0657_),
    .Q(\rf.registers[16][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9498_ (.CLK(clk),
    .D(_0658_),
    .Q(\rf.registers[16][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9499_ (.CLK(clk),
    .D(_0659_),
    .Q(\rf.registers[16][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9500_ (.CLK(clk),
    .D(_0660_),
    .Q(\rf.registers[16][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9501_ (.CLK(clk),
    .D(_0661_),
    .Q(\rf.registers[16][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9502_ (.CLK(clk),
    .D(_0662_),
    .Q(\rf.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9503_ (.CLK(clk),
    .D(_0663_),
    .Q(\rf.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9504_ (.CLK(clk),
    .D(_0664_),
    .Q(\rf.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9505_ (.CLK(clk),
    .D(_0665_),
    .Q(\rf.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9506_ (.CLK(clk),
    .D(_0666_),
    .Q(\rf.registers[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9507_ (.CLK(clk),
    .D(_0667_),
    .Q(\rf.registers[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9508_ (.CLK(clk),
    .D(_0668_),
    .Q(\rf.registers[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9509_ (.CLK(clk),
    .D(_0669_),
    .Q(\rf.registers[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9510_ (.CLK(clk),
    .D(_0670_),
    .Q(\rf.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9511_ (.CLK(clk),
    .D(_0671_),
    .Q(\rf.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9512_ (.CLK(clk),
    .D(_0672_),
    .Q(\rf.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9513_ (.CLK(clk),
    .D(_0673_),
    .Q(\rf.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9514_ (.CLK(clk),
    .D(_0674_),
    .Q(\rf.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9515_ (.CLK(clk),
    .D(_0675_),
    .Q(\rf.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9516_ (.CLK(clk),
    .D(_0676_),
    .Q(\rf.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9517_ (.CLK(clk),
    .D(_0677_),
    .Q(\rf.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9518_ (.CLK(clk),
    .D(_0678_),
    .Q(\rf.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9519_ (.CLK(clk),
    .D(_0679_),
    .Q(\rf.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9520_ (.CLK(clk),
    .D(_0680_),
    .Q(\rf.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9521_ (.CLK(clk),
    .D(_0681_),
    .Q(\rf.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9522_ (.CLK(clk),
    .D(_0682_),
    .Q(\rf.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9523_ (.CLK(clk),
    .D(_0683_),
    .Q(\rf.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9524_ (.CLK(clk),
    .D(_0684_),
    .Q(\rf.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9525_ (.CLK(clk),
    .D(_0685_),
    .Q(\rf.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9526_ (.CLK(clk),
    .D(_0686_),
    .Q(\rf.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9527_ (.CLK(clk),
    .D(_0687_),
    .Q(\rf.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9528_ (.CLK(clk),
    .D(_0688_),
    .Q(\rf.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9529_ (.CLK(clk),
    .D(_0689_),
    .Q(\rf.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9530_ (.CLK(clk),
    .D(_0690_),
    .Q(\rf.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9531_ (.CLK(clk),
    .D(_0691_),
    .Q(\rf.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9532_ (.CLK(clk),
    .D(_0692_),
    .Q(\rf.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9533_ (.CLK(clk),
    .D(_0693_),
    .Q(\rf.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9534_ (.CLK(clk),
    .D(_0694_),
    .Q(\rf.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9535_ (.CLK(clk),
    .D(_0695_),
    .Q(\rf.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9536_ (.CLK(clk),
    .D(_0696_),
    .Q(\rf.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9537_ (.CLK(clk),
    .D(_0697_),
    .Q(\rf.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9538_ (.CLK(clk),
    .D(_0698_),
    .Q(\rf.registers[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9539_ (.CLK(clk),
    .D(_0699_),
    .Q(\rf.registers[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9540_ (.CLK(clk),
    .D(_0700_),
    .Q(\rf.registers[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9541_ (.CLK(clk),
    .D(_0701_),
    .Q(\rf.registers[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9542_ (.CLK(clk),
    .D(_0702_),
    .Q(\rf.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9543_ (.CLK(clk),
    .D(_0703_),
    .Q(\rf.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9544_ (.CLK(clk),
    .D(_0704_),
    .Q(\rf.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9545_ (.CLK(clk),
    .D(_0705_),
    .Q(\rf.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9546_ (.CLK(clk),
    .D(_0706_),
    .Q(\rf.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9547_ (.CLK(clk),
    .D(_0707_),
    .Q(\rf.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9548_ (.CLK(clk),
    .D(_0708_),
    .Q(\rf.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9549_ (.CLK(clk),
    .D(_0709_),
    .Q(\rf.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9550_ (.CLK(clk),
    .D(_0710_),
    .Q(\rf.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9551_ (.CLK(clk),
    .D(_0711_),
    .Q(\rf.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9552_ (.CLK(clk),
    .D(_0712_),
    .Q(\rf.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9553_ (.CLK(clk),
    .D(_0713_),
    .Q(\rf.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9554_ (.CLK(clk),
    .D(_0714_),
    .Q(\rf.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9555_ (.CLK(clk),
    .D(_0715_),
    .Q(\rf.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9556_ (.CLK(clk),
    .D(_0716_),
    .Q(\rf.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9557_ (.CLK(clk),
    .D(_0717_),
    .Q(\rf.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9558_ (.CLK(clk),
    .D(_0718_),
    .Q(\rf.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9559_ (.CLK(clk),
    .D(_0719_),
    .Q(\rf.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _9560_ (.CLK(clk),
    .D(_0720_),
    .Q(\rf.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 _9561_ (.CLK(clk),
    .D(_0721_),
    .Q(\rf.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _9562_ (.CLK(clk),
    .D(_0722_),
    .Q(\rf.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _9563_ (.CLK(clk),
    .D(_0723_),
    .Q(\rf.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 _9564_ (.CLK(clk),
    .D(_0724_),
    .Q(\rf.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 _9565_ (.CLK(clk),
    .D(_0725_),
    .Q(\rf.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _9566_ (.CLK(clk),
    .D(_0726_),
    .Q(\rf.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _9567_ (.CLK(clk),
    .D(_0727_),
    .Q(\rf.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _9568_ (.CLK(clk),
    .D(_0728_),
    .Q(\rf.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _9569_ (.CLK(clk),
    .D(_0729_),
    .Q(\rf.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _9570_ (.CLK(clk),
    .D(_0730_),
    .Q(\rf.registers[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _9571_ (.CLK(clk),
    .D(_0731_),
    .Q(\rf.registers[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _9572_ (.CLK(clk),
    .D(_0732_),
    .Q(\rf.registers[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _9573_ (.CLK(clk),
    .D(_0733_),
    .Q(\rf.registers[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _9574_ (.CLK(clk),
    .D(_0734_),
    .Q(\rf.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _9575_ (.CLK(clk),
    .D(_0735_),
    .Q(\rf.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _9576_ (.CLK(clk),
    .D(_0736_),
    .Q(\rf.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _9577_ (.CLK(clk),
    .D(_0737_),
    .Q(\rf.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _9578_ (.CLK(clk),
    .D(_0738_),
    .Q(\rf.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _9579_ (.CLK(clk),
    .D(_0739_),
    .Q(\rf.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _9580_ (.CLK(clk),
    .D(_0740_),
    .Q(\rf.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _9581_ (.CLK(clk),
    .D(_0741_),
    .Q(\rf.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _9582_ (.CLK(clk),
    .D(_0742_),
    .Q(\rf.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _9583_ (.CLK(clk),
    .D(_0743_),
    .Q(\rf.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _9584_ (.CLK(clk),
    .D(_0744_),
    .Q(\rf.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _9585_ (.CLK(clk),
    .D(_0745_),
    .Q(\rf.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _9586_ (.CLK(clk),
    .D(_0746_),
    .Q(\rf.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _9587_ (.CLK(clk),
    .D(_0747_),
    .Q(\rf.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _9588_ (.CLK(clk),
    .D(_0748_),
    .Q(\rf.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _9589_ (.CLK(clk),
    .D(_0749_),
    .Q(\rf.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _9590_ (.CLK(clk),
    .D(_0750_),
    .Q(\rf.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _9591_ (.CLK(clk),
    .D(_0751_),
    .Q(\rf.registers[10][25] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2821 ();
endmodule
